��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]X	�b4)�Ob��8�O��ȸ�O_�&��*��2����K�I:[�Q�Ar�f=�	 M�i,~4�_F6峹淚'��-So�Z0F:M�&,��k-~�_}������#<	����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P1��r�g����3���o���/�4����np�.1A��06��v����Z��
b�o����n��t1�V*}xZG��g�ǥT����d돢��{���)���v��z�𤸔T�4�,�Dל����ѫ~\��^���9x�6��^�
���4�Lϯ��REz׍��EL�u��;��jQ�wj��:�n��%t�����Y�+	�7���F�Ҫ��D�����Gջ����O���Q�)Gp��B���B�gC+�ys����b���� ni3��:��*���`K0h���(��ش�ksZAA?6?m�a�С���6d�X�)aC(Fn̠ݐ�*�~�����`�"\Ez7�m�K��?��LP0�Y����u�K��;�C2���i~��w��,)㺿t-���5�w�͏���/�|�pe���v�4�<�'|���@�����I�?��[������]~9�e[H���=�U��cy�{��SmN_em״��	�w��Q�%�Á&�!y�k�i�d�H;�h3K~�~!�"߽w\"�}T&�C7?!�� �9����X��,!���`QXq�ς��D���Q#�5i-\��l�=�����H�!����BE�{.<���/���K�rv'*1�{���vorTZX<4�j����ȫ���(�~6�{��OY����"�ؑ���;շa*p|X����2P��H��Wwu��^߭9$����^�*����1$����}^�(C�ɏ01<6�)Q��j�jnSrڋ~��h�%yD���Aս��!�A����4�.�xQ���v�5WSp5$�P�je�4�\8/9�#��I�pK����#Z��
��=��0GB���9�$�;[!r�%�|^�|��ڍ./	0�B�ZF~p)�!ib(��r6D�a�{����?����1'�G*3l�)X���Qg�Idv�OXg�g��n.��y���4�F:f������U�oK�T�7���r-a2�_�ELr��ܔ4g�����5����XF���ɛ*h��[gA�f�t`}}
,e��X��[�(��B�U�ߛ����*�u�EnB�El��]+K�C��D��Jй7ͬ]ĳ�~�1��8��v۩��i`E\�_n|�]���a$�}�u6�AW���� �5��R��A��X&���2��\���;f'G5�(�I���"NtV�Ā�fN?����^�t����(X�j��4��u�O��T+[6&JQ���^��` G2*�y�k�Of]'>�����<5��8��N �vk�����r��2�PϠj�1~D��s��Ж�s��^C�̰�D��H�ϳi�ߩ� .3���dp-��9�\�=�7����/,(EvA���E�s���K�t���0���E�4m ��Lqw�j����,�q�VJ�u���9z(߹We��a���EN���2��r�h��?���B�V�>c3�җ:�$/j|��t�>�ٻP�I<1��G'W�4����r�H���ڏ�'f��#{���܈���`[����U�7��]�Ns<�LWc'��R���*~�u��
;L����K�Ev��k�٠l_(�z���)!�8�pds&P����0+ND<�*O��+	,��a�"2�e5zuTe,Þ	��X��DJ})Gk�Tױ�yw[��ߙ֓�]��Ĳϊ�w��C��M
F�6�E�b�t#��kxù��C�]���i: xtʍ��ҐM�����:�I��J;m}H�1�58�uJ�9F'$$�����OK����X&���.ק�{a�/x�jr(AZ2�:p��-�:�M\$-���U�15��Zؘ�����3��u��&�;7��A����<]�F 	 Cv��D���Ʃ�W��Zyk���Oh�Ug�	f�c�&��f8H���A@J����ƾM�̅0_܌��v%ʅ�P���9�Ւ_t����kW�'��V�BT>��(�/̼H��w��o!�*�3|[����-�֒n��|�aD3IMy*7}S7��Z�9o�
8>9�3���������F��^�f�i�����(��V��*��/�AkU�4�i������/�'���ܦ��N�|{���̊�"�h� Ӟ�E9���>�����C*½�+D{	��I�C$`�zE���|�a7����T!������u�Li�Eӧc] Njѿ| }R��
(���Рc[�P����~i��	��3)����p�.i�A��.��-n-|�Xӆ�����U✗F�Kvӣ��0^�h�V �ǰ@��P�o���J�������b*7x����TÎ��y�i b���J�邁��G||5���4�C6���3�uGZ���?| �7�p0�#g�7D��PY�i���*�]���E�;����nGH�lҥ�	T?�ؔ�,���+�cgO*F'����:���=���E�����l��W��9e��`��>f�r\�"�D�U1�5
�z`�ф~P�J�ЦzF(� �p7��������DKM�5��y'	�����{;�=Ƹ��naG�d�Bs0�RC�eӪX�̄��9 �I9�	���;�8!'���0��X�D�O��{҈ra�՜DJ��|cZQT����z��z�ڑ�<&��uM��iU�;�,Lt;��X��ƥ�����^$���?���.��(Ȉ��SSZ	�+�ՙs�3µG"w֬����������8��ۤ c�������y�X���y3���ynUA�]Hy���..��c_W5����<�x�zL�\AT�q���}���_�=� �р}0cE�hk��/��up��@�ņ~�W5�����3R4"��Nh�����6o�,y~�)m��-!Ĩ�H�ܕ[���j��ˋ
�?p��b-Z|�0+��t�[��I�"�($OU�b̀-ѝ�yF�ѫ@[n9�чrP�$��D���F=��̬��Q�ǌw�C�p9 u�;\�x��nCt��ms|�pšlz�-��3�?P�Ey-�>�^�Ϙ;��/w�p i�k�����W��5s��t���?w�YS��U.�-oe� /Q&pbX��\e�y�$z��Q�v�VB���N+���~�Z�P��-��=`��p%`��<�04��~?;����8��T��|Nr���S�Z
��@��t��{U�IK�6;bR[�7�w��A�Aμڌ�s+V�ڙY�G�����s���D��S��
]�����B��d�Kʰr;�7ב��*�����,���0�f��8��̺���^�Au+5����*�լ�������ŵM���v� W ï|�EO���Ʀ��z���W��@��ߴ�����F���S/y�s.�>�+�"q�0ũv��T���־�ґ9�m��ߓL1��'�c��"�1�Ɩ�-����{�	�A4e�m��i��b�� ��L7��~��%�h/�eL|`��ٕ�G���G w�-S�?����[��m�?�MC���E4V�p0��g�d�r��L�.p3�M��?q�Q���������-�b��<3(壊2�Z]ߙ��ȩIA��
a�Q@Ň�C����=8���b�O��\̼>>~�'϶!�ʾK�f�o��q�ߊ4�q1�V4./�m��$2�N�ۮ��Ô�53�wIe��#]���FU���+գ�f��
���)b[�H����l�N�hx�|�����u	�\��� �qN����n�H�����@�߇��Z��g�Oݭ���2�L5�He$�.�����Q̍�Ⱦ(�Y�3��/'nE�Z/�+�s�
�Ԛ�@����{���QB�L����]��ē�}�^}���9 β�htE��mJ�L�T�j��t���>ӽ�q�-w���?�X-���v���ج���x/9^T����:m�4�b�|"�VL>d'dR�z9PD��C�.hfE/�>����"zg�_,?�[��i��T�_+v0jLf
���Ō��E5J��O�>6�vS0��apZ�8���B�ՙ��2dsrCj�����K4�ay{Dv�Q�Ud9N�����*'D5��t^�T� �Y��G𨄹�V�T	�wm��:MT܈I��tG\�o��S�[1�Q���z�BӀӹ�C`�����(��uQ��ڀK��Tf�J�;N�;8� C�ӈ	�y��mz�HƯ=����)�@��&P'���o��zR��X-��.qW4���ų�ڌ�i���W&W�A�ŝ:�w�Ӈ] ,��	�Q�v��ϧ1��;(z�H�t�x���ĵ��L���m�(AO�T�;r����]��Tdo_?x]�_�*��G�i�� T8�1�jt[CcKHc�ňn��Z1;b����%�^/��t�<�A��FJ�_�����9�̀Ӻ�ļQ.�r(*,��=+��Y��ܵ>�cbT� �;�zF�8������L�rm{5���C��U��f�����5�Y�W��T����h��	�jF�[�-J V/��z�a~�%����J�H�풦�PWC��V�C.�ݦ��3����~����nN��Sl)idAI�"C���"?���5\��p����e>)e$a�+E3{򹆩�hn���w~K����aO�Y�������2'u�,5�kI��Ge��P�?G1�}#U�D�b�{Bw�W=^����s�հ���ߏ�j����� ���A��S�x�t6~��z2�T����峕��3�l���|:>n*�;�-%s�����b��t�W���ɠj�+�1c�ZM�c���˥2�l��{�T�`��My��a����"�~�gݽ�Le�MG7�?��!D[
�af����QFx�TjyF�m�A U��G(Q�#~���,��;ǈ�wO�ьؒk̃��[�E �
w +��u�oK��K����N���j�4e�v�p��t�彜���/�]�"��'C7q&�{ܝ����:��c���4C�)���x�����b���'���6�kD�]/�l�&�\J�֧ͺ=?%N�j,m��x��jְ6��ҷ���1Z�^�����lnD�CГ.�h���$I��"��$(=��P�d+�M�dTb�:�F����׻X��������}.\
8�IQe�p��6m��<��ٞS��x�I:��E@U��w��X���!+�!�W�k�s!XPѲ�,��q:2&�Mq�h��~8�0�0��q�w#N)Hj���ޚ���*��[M�,S��X���R��H%��j�jN�*!�U�M*Xb�Ҕ�e1�w�ҳo��1s7�k��f�W~_ǟ���m�8wJ1ȳr�Z��{~��(%�r!�a���hӖK>c?��?戇fG�C���y˕���~o Ծ�I��2���F�G�OK>�~w��M��7D�RK���|rU�,��ΰ�՘���B��ڮ~�euq�5�����C�Xĝx�M��^;&d���Ç�����P8�#�\�o{"AִT�쾂X���z�a��#���̝(3��=Z�=JՎ�'�a���K�d���v��{#���ye��x;-�j�=o1�|��d
�.b_�����i�N�nF-?��Uz�#����n^8yi�Z6Q͡G���ˢ��=@�b�H
�W�����Ɋ=)�	v��Dz6�2�/��O�^�(��� 6|h� �G��S��nv5���Ԝ������Ti�&�t%5b�*� ��
�X\5C�t�Mɻ�"w%k�����櫿�`'���W1f,�a�����3�JW�)3�_�(HKL��g�gh�[�s<�8�i�mH��ɸ�t4E}Y��FyO s<�'d�6D�0w�S6��z�ʿ��5̠����p�J����u��	��4�i�j����,
R7b`�<^����+���'��\�{��	>13Q�|L��0�[�3�T�����Z��V%����t�h%8��*s7��#���S��W6�z+D�����򒌉5�u�J�TF��˒�;�S��K��*�w����OR�*�WX#1.��!�,݆{+��ُ�?���[��P^V�f��֚.M��1�b�|�Q|�u��K�iC���G_-����`��gH�{�{��s4ˌ��z�u��dC�L�U���+A�#�I��_e�,�p��$*���OF�7=�>)�?/*�^
��B:T�l,�:����rM
�>��7���'� ܥ�v�zXU����9�[�}���l����ԸGL$��o�"y�|!{6�(��e5�!;�>�{�`�){��R�5���$��'�kc�@{y�$* ��x��h_��I)}��>�/?�_����R�Xx�W[�Y�-���}�.qf� �H�To�C�93]Jß�:uL�!�Z���e!�Tu͊:8�Ѧ?�gc�/�S�8��ά��T��2(V�/ C8�y�������ڤ���i�����+͖��p#��~2��Y �h�R�6A+t� �Z�n�ť��#R�Ho�k�E�k��qy��֌���Ƃl�2$d�q��Z���d
���5��$F,�-��0%P���P.3,��LIb
�E�rlx�L
�f����:p#32�6$R�U�����n�0.N'��u�O�_�Oy }�<n��R�����[ax�EA��J�.ʦ�%�d�Ⱥ_0���+�h�b	2O�G'#�� ��p�'2eČ���7��o�Dt������N�e��w<�����k9��Xܓ�;�F�#Օ�W���Z涗5��
���cxr'�L
|�a� .�9楦@=�N�F�%�3Q���uio��:k�䨫��!pL˯H�훐�W�����_������(�����T@��*as�
-A�g� �]^zB�R*1Y~��[�����__�xɴ�>3'��J��yl��!��\ɕKDu����;|�����Wu�+� �=G��CD��oZxo�z��c�e�� m;F �m=�* ��n���a�l�A�����oZ`z%=��6JZ��*&�j�i@��U��R�f���'��	:rˈx֘�%"E���"���rhs�ϲ��H[�P'��)�!\ �:6h�n�h:�O��� ��T�ZC�٩�
|��k���S�a����Y��#V�*���X��d�7)�Gv�96�� ]�8tjm�7�:[��<1�{b�7^��E� �=�'�_/�����\KOx�tȿn��1��A��K�Mn$dVq]�63 ��-���B�T j�LW�-��{B@(s&�����AymawtgL���x}#��JL��!S�����)�g����&@	�[�5��1�������������g˶f��GqM���hyI��$���JT
�<E5�l�j���X�DC��	L�J\��{���m=��[��yAb��躬A�Uc���8	ͨu����2:jH��ѥg�a�F8�G�`�Ul����c�0Ø�M��'ѡqC7�x9��"�3o���FZlqV��+L����"��jsH�7���C���ΜP��j��F�\r5�6B*��^��	V���e��__R}�.׈�t�WCt?���?PM�K5("c/��-g>bH+��_�H	u�z`�=�c��*�2S��^Y�onJ�3��}K��k�RH���1+k,��`)l�]_D���z���5o-��f���c��MM��x,�X0Qb�a�A���
�`�Ã%�C�Ah ��ʉ������]�����Jl]bF�s�eߞ3}��,��Z���>dH�ǜ���"0�LrC�	��FJй��>]|�vÜ�k��}�Os�����.��N-{z`m�)i�z)½� ���t�'3��*¥s�N_ ����ܒ���f:*V/��ֻ�d"j�H7󂐑�0f0�Q1��n�$B��u_\#i+���~S�K�@J2/6�.r�u�.�+/�b�t<��ϓn�q@�9~9?S���c�t�I'0�����ǎ�����kƱ�u�;��b��j�g%T�?�%�i t}+�d����G��Y�e���S��O袜�1n�ﲱ�FD�p?Η������zyP7<8�hF�/��+�
{_~>��������M��Xʀ�^�������7�:B�A������<o�7�	�"��e.~��Mۦ����C�PY�O��v;A��b0�/_B�_ݾ=��t�&?�ѝe��Ǩ�,3j����&��Qg��ؾ��H�,z�N;~��w���R&�*r�/;��X�00�V�o�Uډ��m���W�U]j/��R�w ��N�2Xod�o��s1����B��B�@Ą��� b\c�=�<�O��#�N��ar�Ѻ>jV^�1X�rJ��շ���x�c7��'ҋK��AT�����Z� \�"b�ƣ�!�	��**@&�G����r�dsf<��L�r�}��s���w�RZ�vvir�6��q���}ɥ�������T�d���>�:ϗFS�J�������+] Z[`�����Cd�B�Up�m_P&+%q�Sո��d����㙕��@#��̶�>��n#0���}��s��]��������pթ��E��a������S�7)����v�~Q䛵���{���z��쟧���$Q8ٸ�<�����7���8�ތ�[��*�Ai!S�*[mCȷ�JN%}��3��`�U̺��IZߥYlS�˦�K'��+\����T;��ȣ��)]?�Ȱ�[���r��V>�OPR؞/4эqL���׻u��b�L�<�M�gP������4�ފ�W��%�e�R5�����f�R���F�B�Q�a���M�(v&F>i��ݦsr�n�	L��2lb[8��q�����u>%�k����H�5!.L1�&�֓�})��9O��|zh�aXV^��=���(ުQfU�Þ�jK#��2�U��MK3�Ɍ���p�^dCQ5H�+��ӓ��-3���2�$�D!�Z��#�p5�5eq�$΃Až��V�N��2�-����B���]�uҶj|�t�d�����JjB�m{vA�UW0,�N�_M��)��h���h@�#���{r֕tm#�e)A��@C]@I���u�+��������{q����!��V��M��\CѲa>�+6w;&�s���}_�4��S����>��o�/{�^z�dV�b����e~�&@m�3�~l�ul���#�<�&�kWؤ�ek&C}�� :��w�#��K��$㨧2mSn���lK�=O��MgՌ���f5=K`<�!�Ebz����`��dr����I
��[ꞃ���lUU��?��&�ٝ�ʷ�'2X�٤�(p� c�G�wg8˽q;Z�PQWD^|���&ԨW�Z�;e���'�2g=\S�n1L�g�m�ECҿ���F��4� ����xt ��"�nD歳!=�G
#�p\��X2�(4�=#zR�.�<$��/��;�ټ%Y��܈w���'V���Y�P�O#�o��0\j0C�;�5Ѣu�0O	����`��+�b����-Y�Z4H
"}+B^H�];>�"ʆ@�ץl��*��ւ9�T�����Ώ��� �9GŊ����w��l��6�wuDr����c������UXg�T�eϛU�� 0F�
�P�j^��q���p����˥!��
�M#���ЮĊ�����"t�������y��$>F){kT����e��Q��ݜ����p23��#c�c�yB�Ds�	'���܋~�J^Ӈ%���jj�UPn��� �yw��C�TQ��S�A_&+B����;u��-��Κ� �[��ʚ��:�8��x�����x�
 �8���@$���h��Yt�˯Z6+�iä�䑜=h$I�������h,�E�P'C+�S��]���Z��IL��!"NfJPy�}�+Zkn�i��tkP�x-J���_�ի�	�椚<��FΑW�0����S$�ҳ���TaxP�^%^�7	�F�d[�X=m�c*EL�r��w,b�U0�eP�����j�`�Q��]*�ͮ=��%l�<!�
��0���S�
�t&q>C�$U�b��3w��<��:@��j�rH��a��Zª"�.�c!�nd���m�����n���Cs\C���`_CІWP�)�h�$���ҕ�:F�Ѥ��x��U�9������"h��Z7a�q9s�0��fC\{���9�z��l uRt��J?Λi`h��q1�����K��F���N#ߡ��O?�jSxӰR�q��b������>�,��S���Aǚ��Q6��l󩁫$n̜��꾐8�ld�&#�`0�or��;����j}ķ�K�eO�lu�@��jp3�k`��xd[G�%G���4`mi@+�Τ|��\h&�_?@�k���p\�e;:�o�-63.~�yA&/�.��U�x
�,�+�¡�����zB�e�����G��"v�v�_N��!�1�<㭜��j�Z�ق=�IE����b<�͏�v�Z��V���v#�܊ُ�JB�ֻ<�̨���)P���؉>9{�*̘#���~���)����V�`~�F�o�nݔ�]�����/鑿�&s�&��K�Bd9��tm�����
��E�z�0����0>�A��aPX��Ӡ���w/������6H�X[��)4�S���8Ꝗ�[E���]���G�}����4��U�i�ۂO�~,Y��~��&�3z�/J�"�q��y�gDXߕ�U(�?��9���R�v��e��Ł(!�?�E�I�z�j�$�A�d܋1��[{��[�����_u�29�~RͫA�R��J��۵����AZPo�㬒W��^�u�Q=_1 j�ȳ��Ԏ�.z����Қ9oI7�R4������f3J��y.I.�Pܞl�u�z1������h��B۪�P"�����M�b2<��rQ��N*	�EuQ�<�ڕ�R_�U8��p�4�����|��Co�m�Nc�m���\��U�o��c���?J�l�ZQ!llc��-�z��=r�����5�����I�v����6 �V�aa��M��҆����t�*m�P=!Du$Á^{�"q5?KҒlZ�l}��>p����<t���܈�AQg�s�n��p�(/�'��IZF�-�o4��y��\9��Wm�ϫTF��#kt�=�ؓ�h��b�?˟���A��S�Ts��q%�	���*s��λ�d��UY0ة�Y�=�;�|��<W�5k�f��qekL�^&�$s�7��7hr�X��?��	�q�X�=��mK��t�4�L�3(���	5U��͌ȖwY�d+
�p;��NS����6e��Tv�dƘ3j�l��3%��T��9����h�E��M�=�H��/ݸ�����ge�=�(�ӊ7��چ��U�^���Y��N�=F~�?��=����l�k8�g+:n�&^��|T}����W�g�_��g���8RI�si[A��}d�T-��_5C��L����"��m���#r�N8C��������:~L��"�g÷^(���/LRV�=S"`M��r��C��kR��\�="���O�]n^�G=t滣�4N�s-k�Dr�Yˑ�:T��R>��R@����Z-p��W��Gv`K��A�阤[:���9�9v���L�����Y;�B�3(y�[a��V�.�)̉��<ru�aVV;��2�Po��(�A "a��̯\-QN�����Q�����p��Wg�j�[��������R�[K`@�$o�Q��~s9%����0ʂqfk�p�{�h&�~:[	P�1��W4u��f$'�3�Wp��_NF\{�LB����~-�~�ۓ��cZ�$*\�����ʃ��l�
������K��#� #)��3�����o;�4J���=�:PY��S7�!FI�@��3�nl��1ǆ�.�G��u�8�hb9.!����Kr9/mE�[�Y�n1"4N�FTK��-]��[>�  �\�b�o��-��#�5%��$?�1�1�<ak���3Z�ס�W�.d�5�}��*��^?~�MAJ$�Ϊ�@�ԙ-+ �L2z��`��܃���_~h�߻`<�"ndR BJC����,�t^N[��tȾ���)
�f���V�qB��'����f��9�#0��O�AA�tN",Ʀ5��w�g~�����~|z�ȉ6D�n�N�
�(k]�jp+^C�{���'��܂�dV�x���mU��m$3�
���؊i����j�eOX�Ӕ��̓*����{�5gɫ !�Y%(�h����.��@�$t�y2�:͘A�S�;�X�[�34:, xK�����;�	fJ�}EM���'�+Hj2�m�e��
�}Ph: ��&�4B����s� ��.�M��=g)����kY�ʊ> ����C-V������+(���D��
>�o��&S�;��
|M�ѻ쐚�����u�r�4>Ŏ!8	��|!�ǽOF��?|�K����hދ�o6.�ß����g;D��`�e]�v��x����͗,S�Ȋ�`�׃�^�%����\&\'#�*���_��[<(��ӷ�%�5a{A�<s������R����s�yR��C�)<���ݸΟ�^g ����FyUN�]�Z-1eʢt��C������*e�'TH�;�7�\�[U��׻��Y���Y\1���W��t@��/s�)�t󘳼8��>�7�n-�I �N�P�ɈIIu�׷^�k�N��l��b�P0�P;��1���r�~r7��!ȣ��/pI����	�9�0� 5��g���� M�F�ކ�t��.w���n��s��A��f�c����=��&ɃI.5 )�w �HSH]��V{�,��3���<%�R���,'{��</��z��"A��1�G�*c菰)�3�]X�p��W�����\�Y���8�}���2fn�0ڋ� ���^��]�3���t�{��,���޶��g�a X��K��>��oV/d2�����)��JA?X��g.��	�+n�y�4����>�̣��d�.״2>�Z�KCM���s������z�o��C���-�{
j���=���G���"X��UH$�@u��Hw��udF�F�Ƃ������!��s?���L��ǲ2�B!sy��-�{F�aJ������N��&]�X��(9�H����Qqv���"�<��Q~V����<�Ph'���||l�A3k ��"G�������<�5�Α�	_V�`���-��1E{�g����5)a4�Xe���S�]�TSu�I05�h��b���,�i����u�����Xj�v��K}��G��O&յڐf����gu�E
3霡-�k=${�2KL�jc-dbk'c�)?���$��A�R�v:�_�Lx�χ�}ޗ��b����F�Z������YZ@�q�nDe�{��D
��x�$����'3�C��>�-�I;��90�6�UK��H���ǜ��8q8m�J6��A)�`Sy#�F��\�;ӇvHp�-AҚ�L6sO�����A�l��~�Z���U��pwst�����H�㽦����Z�+ϝ,�K%�� ���d�,\�^M���I`,�+.���'5�jG�\՗#6
ĒI�Θ��,��ʙ��,:�@�y!ǔ�c��O���Q�r�v?�hG3������C��2n����m�:w9��7t�$�t僌{8��]�4�s��"��6�����2�WX]Lpk�NG^8W=�!�]W�te_��E�8�g�֮ XJ2���/�,�Ī�F�_P�ŵ��K��]�jp�8�_�_%O��n�P0-�A�.>IEN9�[u�t�
v}�� �=9��LG��O<��"�Ay������ǠLd"��|5h���Fo<�����V�>���'�Ӕ�v���=8g����`i��3��ǌ���Y�,E!�~�y���ذ��G-��6;��OhC�WXf/��Qlo���^�2��A~2�@x��a��DWFcdy-���˜�ɀ�.����+07���r���ms���>x �ݨ�k�/%����>�_ONPw8t�<r��a����"&_3�m���UR��G�V�МO�F���o�nLă����j`�nl' oP��f"��>����"p\[����S�&�H6cY^:�r?��dҁ�E|��Z��~���뙡���7��(}��˿AE�\�6�u迗U����v�g��n�㥧e��-��J8�/if�����~��Ie�F��.����mZ7�9����d/��́m�z~�t��5p愓)�t����i�� �Jh$TMҤ[E|���������3�u���O��y����`xTra��"v!|��Q�Y���nunQ�ޥQ��a:kP��
хi���zL��YĲ���&/� \r6���Xc����?�m���b���$K!H�K?�2�i��(E�=�������5�����_O;��>��PZ����O�c��}G^����1Ӯp��2�b'��U{ZL�MZ�I[#[��9ݙ5�U��������3�"]&� F�&��9JþC^���&����$�U2��x���}`ӖlO��,���E��r��jjߗ���
��%.�\��+J����:OT�2xs*c�LEG�Hh�C���3�ň���g�O�c�l�OA���o����9~�i ��b��,!D=��qӖ����B9b'�.�#O����?�gkZ���7\@3Ym�V���Jz�H���h/\�3�l��<@�A��VX�R���������F���]IJ�|�悎wpuoS�ܹH[(A�ERv�Hu��BG{�}�`��[�0#�I;�2�3��g%���3J����Pw�Z��HPX���=������H�Q+�`���B9ˆ��.z����6�J���uQ����.*,��綢gA��<z�{��ύ����z�.Sux�ũ���z��/8)�Tg�L�\���'pmϽ{cD�l���!����uybj�����.���T��%�:��a��f.e���T�AS�H֝n5�ӑ�Z�l�k�#q�3H/�+��9%H:�l�U�XP9��`�R��~[.T4Ē�Ե0~�ǒ=z�2}��dվ�M;�ed���4W~x��sû�,u϶d�����qE�Kj�c����?i�;�Z�!�r��_�g,8D���Kr3=v��؟r~k~\b^�ꐢ�=�
���FFK}��J�[��ph/�s�+��й-����Z�+��|���(�?�::dN���,����<�4֚�9�# ��ˤ��v�IZ�;�醾�9�ͼ�.�{ך���(,6�#I����u�t�H���-,���u�N�����߮~�:
�
2�/�E_gHh��y�ǀ~ץ'��.ǣd�N�j��&U�T���T�z��F��$�,�<��K��Yt3����&�Y�n���x[����6���@�� ��M15��������Pwr��Ù�E�<�2e���!�{�'��t����59��#�ԏP�W���Ck��!M�0��M]��}�L��-.������c����ݦ�,�y(�5mEe ���ŊC���vP~<قc�/+�Og��?��f%�b�Y���H��üV6ah�<�I*�a\�y�p.�E3l֑)��T<��>CװE����G
Ƈ.���&zn@�c�0���M#�~�j��2Q�P�� !��bn��x��_4mC?y���羣�����9���y��g����sRv>�g;����,�E�ړ0m�(����m��z �}[���-������5�RҚ�D���h����r�<�Q�_�i\�R_�!=Q��@��K�4�:������3C&*":84ԛ��n]�O�%��v3�̅��y���8äD��`i�P�-�9;4[0�,nRi>�_��'5�N}�m"��O+�)yt�Y��GVN>*�Vf%���rK������|��,S=]�0x��ŕR'$Cᯍz��#W\��,�)4���Y��}���}����;劮�$��,�S��H�jP9U��A:�r�E>r��ʲo�y��]�b�~�q�-�ǇZJ�}�N	o ÎXa�l�d�Ⱦ:���0q�lj������+��.�t��l��	���T�k]�^��'[��Ϻ��@l�'��)�����*/=��4H�Y���|���}�b[ˊ/����KuO\�j����4��6��^�\����6*�!3k+�$�@��H&��d�!���r#7�Uh�0_5�e[,��s���Z�F����1�p�6����=�
0�Y3������`�PݬxS/i�'�;��|�fry($<�csH�E���L��ِ���%X\�8��7o���t���׭7x7�H���͂�u{3G�/؜��G����T�&�D�A�5�	��x�!E����qI2jq`Hy��P���Q��a[��X' ���N�?.`b#���պPG��NÅ�%X���o������b�5D�^۴@�!�.�t��bH�F�[��Bq|�I�?~������i���L�`�r�K��_���O���-X������i������s��s!���L�����\a�7w��K3(��d��)��fE�����2��S�-�oDSCo������o�o�6������qU��R�|j����.�j���^{j/rZ$�Tx��Gr�y»�IAb`�g��8P3ʛJ���yS4�G\\,�Aj���N����a��Y��@�R9U2�b}t�b���q3`5��4��� ��m�<g�R����c4�z2��	0����枤g�gS{�J\��a#"l~�E�BN/��rEw#-q��� �f1����~*]%	��Q�wJf���\И�R�tdYA�D���-�ryXfU3J$�,�+��\(t޳-�� n���;��.殯�c�-��������J�< Ы  B���7C���5xU��(�v��D�l�)N�@A^��g�\Ջ�ȠF_��p7�g�S��P�'�@��9�S��ft_I��p6�g1�8n >�h2�o�!*Ysw�7��7?�(�w z6�*%E��^�U��-��e�3�h�!c��J#uG��+ 9�R�=���XQ`GȈlJd�j�i.���ކ���$=OY��%���ߌ�C'j����̲��KU!Ǔ	���.�xv1����g�ylF��h/#͐c˹�/M��y�b��!.��oi��@�H0Xv��S%�:~k���Q:�&߻�m�"�D�%��޳��*�)�Y�[\��~Y��e�:5���x�V����;�[6	"8<�gO���/R�1P��p���@|Odg!�T�R
",���Kau�|&!k�r$�5~�'��ڀ��<����U6���Y���L���h��q�MK�3�����i�k�'��+v�6Ï��N��J�nR�JV���;o��(�~������e�D����>�5��:R��2aΧ�����t[��	 �1|�S�|M�q���F�p���i�~�St��-"�p%����p�����r �eb�;K#*M�����Q�$@��/hB���H@��(��X
� rN��X�[�80�sY*Z���	йL7r�6��F۱&�-p'5dˮa�;��A�~�2DI/A��~dl����I��{ou�ݯ�Uz�T��^[逖8���IE�N��-�a9�5��I��l��p	i��W�����x�`-�·N��iJ�����Ys��z[����l���_
�Q��:H�4��N̗>���+�֪�+��Oa�<G]�X�?�A-��5��e%#x�e��*0���@(�E�"g�m�IFq�t֐eL�����Ӈ���J��OrU�ϒ�$���~�CWymY��B'��rd�����m5&Ag<��D�^����\��<�t��e�8BN�C��B��WO��U�1��&'7�iL���֕#�&[�;��5S��ȼ�Z:V>/ �Na���}¸5���hp�\�����P�K�Z���F����9b�މD��@� ���%�L��&�]�m9j� ,?��G�o������S���s����vO�`m4C s�g�����c�Y�Y֭b���0���u����_f��`x��'�/�(-�*+#I�3E�/���3;�ge$g�uC>�s�e)�I|Y�i�4��T�Y4����][�^�؎~k��f�Q��H�<؍���ɗ�j�36�t��(�К����e�^�L|Y�9��0�h�^��?���wy�j[/�ݵ:�?L_9���
Ԙȗ1b��]d�ױ0�@7����T��u��mX���Ƙ�qt�>kѥ�)����ӣ��!K�)�뵚�t�L��f���nV��~�&����ל1؞�r.r6X��K�gP�$�{Xk�# �:��=~z+�?�Yа�����gƕ�6�9�X� c( �e�R�+jl�<����d6"���E2��d��֟��e�/H2oAC���EL���ڂk��O&B�J3+�����kFs]����[���M��1j���4�I!�ħ�W�K��c���p�qc�h���������0�YT�H��}{V!ˋmK絪f6�+��h�o����v�RV$��F`j��^�2�_�S>�9�$/z��wSJ)�u��=�qn�d�MmJd�^S�
��9(��W��1�叜�D�ɳj�q�z��������t����d�ӜǮi�,���u��b|o`6�90E��H��q1�5 �(��	����4����((Wgw� JzU��A9����C�$�-���O� �0���V�l�.1�M�R�e��b}�"���_�};%�T���>TVū���/�z& ������ǉq?�ZX��F����{?0d5�N�y�	.1k��)��ܛ��9�[����X�"G�Ɠ�h�S�Dwq�
�!eŀ=ǢC�x�c�9c��u�+��h_ ���E�^��g �J޽�'G?R�>����!1\��]~���}E0N����~y�󷝕�[%(�ܠE�O�7r��v4TzF㈋�C��p�hϕ������6k���?rD�_fi�[��
Qx�WR���X),*1�p��qΛ��3�b���dX�9L�����P��!�q��:r�%\U0�T����j!�B�j�7*}��B�9�Rm+��2ٚ�r�p���@�R�����A&7
%��Zz��4Z�e`ff�0�����B�`�M�����E�}Ė��M�sw��xy.�$I�Y-������Ԗ�=<ɻ9������I����o�ߖ8��t�Q�k��!���cf�;qw�a玄�YZK��fVQEL������ ��#��Ow����u��"���`��#���&U��؞���>����/�⭥�[��d�k�v���e4+f~��'?�C�~]�<��'�����\ƶ�m0��a���|v��· �t��J��՘	D�Z����]E8��I>��Rh�[r"�������W��KG���莒��9�$Ϣ���7Sk�1�1�upJr�3+u;���j;J������حJ��Q��MC�pj�f�6�������[N��.�P��!N����W���Y4p$�=A�W��=�S)Fk�r��sJ�Kϓ���\��}�g��s�K�k�ng_լ��D>��f�rb�D����wh4�z]��!��]��S�0���s�/l����3��׉p\�r V2̸�UU���E����>�5:A�~�]������) �´[j������ۨ�-�mmo�w i�/?���)�k|�.M��<�eň7���i�g6CY)ҋ!���H���ޫr���<Ⅼ��z�y]9��Nɯ!g T��JYlX�˗o�^������T!�yN XgZ𔕵�A���A7/���|:c<���G�H�3�Ce�����d����]ɧW�� ������l���+2�j�������Ս���S��e9�԰�11'+stL��K��Dڿ�����N�ao��i�ג�t�QE���{y� �fe�Z����q:�z�ԙf��AV:>�R�mI<A`�)��#q"���a�W��m���Z+~S=4]?�3�?��%e=�����+cm2�����[?��� �C_���uWL!2?Jj!E��Ac����8�Q��	`���� Q�}Ӝ3(z�,5F~r�Wp_�v\�!��(ڎ���{�H~�-�jv+3�?�˕;ʦ>���k��H��(il��^�ˆ�r�z���16�����T��/� TijTT��c�6�Q�k�^��bxb�G������j�C�.\�E�sP��&�ݨ������a�'4����-������7x]�ˬ'��+M��Cpk�^����7�;X�o`�m��F.{�(��G��w�DQ����
D�fXeS��I�Os	���E-���``�-��4jq|w�^dڂ�J��X �w��x�Za����`$SA�\|������:��ot?f�y�$۽&,1_�Zg!i�オ��|��Ze��)����E�h�T �ab�̟#9�4�_~������M�E LF<�)V{�{��.X
)��y��W��cEf*�̼ǟo��i����������7�(^��1���`FC ���8���=�?�����M�v��U�/&�C��!^�F��B123�-[U֔�#��= @ev���GXh�����{D�B�0����>�֎K�Wl#-aZ� ާ�h���7�,o7`��G����o���V>��t�3"����]�[�2��5zT9�ѫ����j��oҋ��GX�HϠ�;]y|�ԏ�-OznH��12�h����(}`E�Cx���F�綩��.�.��#97��Q�&�;��:���U�[���H^�(gJ��<�A:6�h�N�h�
�w���v~���ڭP���H���\������d�:���@_�A�硿�Ύx��zU��q"A>$�Ј�r?����n��Hʆ��S�v �Jc�ǁY4E?�\��b�#m�k;^�e7�p�q~�q2w�>~�0�2��?�p�M���(Y�R��ڝl�*�������k�����{Sr)5�5�0�w��Uy�J�ui��Q뼿{�.��y;�ص���P|�����~7����OBjr��!j.G��σ��{w�k|d���4��kp�~">ˀ ��]���\t;��"w�F��Nc� ��z�5V��ɗ�+;��I_R��j�]���"�)�߄'��ӴOd1������B:Y;ڻ�-)���!�}���X�2��+ 	��;튣�N>��p�ͣW�*bk0����S��?{e�bѾ=]��6���/�F;��d������F��~�3���p�0�XI2�������$-K[��u�O�seP����X/Ο�=@kwx��3�0Y�.;e<t}�J�!0Ð��Ღ	~�8����F%V�4휲wF ��;�}����a��YY�"��͚ԉQ�2�s��l
(��z��ht�Uiɏ�Yݠ0��aR�)��&��L+;ȿz�XT(�Y!���UEĐ�֖�{G�1��8�A'�l.i� E.B\ɂ��K�r�GI���e�e�1�#*�3�ȚŜ��3�ԲpV?���A�5:���&�` �ju����?;ʙh�WC�̐��z�����u������6$�٫!H ���B���b�7I�V6�O�6�9G�p�@�d{3u�Ƕs�x�-e���OB���G��(����l-�d�P	6G��ω����"�5	� P󴃧7�܀�N���dx}$�k���ޣP"~�X��wGM����"��>��F�^Ω�n<QGg��T��ٍ�]�˷Iq8�͐�4��'�ɏ[��k�l�F®��B�~/\�U�FZ�7�8��1��)�g	�v�L���UG̿��d����s<C蒲1=�A:2�(�Ak����բ֔H#�t|�M��5�?���u���q��M|�ǖ�('����.�d��m ��O����g2��.c�e�/���I��%�VLcD�:��\���$��xI��?���n%�����g-Ppu�gu%�,NIP��bD�5a����9ߊ7:W�⛚!v	�JBƶ<�<���͜o�mdy��vAխ��t�=.W��S�=���=h����aW�Ԇ������IX�I�j�c�-F �dO<Ԡx�*;�2������v�����V ׷�͈�x�+s*���A��oЛ�&SN�=�M�̮؍"��'�Ӄ
s߿�2��1�;!�BS�+u>��z��*��4A� +'o��Ƨč�KƵ��l�h1���? ��V��*�H�I
���Vc��v1��n��e �cp���lȪ#�	m�22��*��q�Y�kH�N;2��]�.4����T�������/#���礢�2���rKm���i��i)�(0���ʡTͻ�F�<jYhr����2�#�^������Y�$�����k�.%����\L�O��;OV��������=��^��с���
�Ɖ�qM6z�rh�`��XW����=u�E�q��3o�V��GtK��	����~�E^��䕋�3�!�r{�꼯 A�pD�.��d���\���&~��z�q~��;=8V�*�R=�f�b�JO�ڱ
H�|�u�a۶��V:�61�t�J��t�U�$'Q���ώ;'���i������Ѫ��Wj�֐�{��G�W�1Ism���ͼ�~i -��U<�
��o��GR�&���t�/��w����e��Mv���H��c,��3}���ш�s����<����(�3���5c8�3?y	k�����2��[ST�b���Ln�&dp�í[V���ej��ȴ���q���v���	�es]}���xop���"�����m���̔os�0��C*��Q	�4��;v�=�f0<�1NN��|���p��G�5�n�Ѹe�7�ڭ�F�}����[���~^��Ϛ);=D�Hd.��&��^���O�E����I��\$��M����\I*���h�w�p�`En �Ƌ�]=�6L��&�r����G ���/S?W�2�f^�Æ�n�07��en뷆1b�pg�y>�H2��iH�}���?$�QR6��>��Z��ɵ�����kf"	ֶ�Bc�'��m�Ϸ�D|�2�!�y��5����1v����dg�а�����S�u��A���Лҩs�F(�9|�dOy����H\l�h̙���1�0^.��E�}UYq�'�^D�O�R~F�;\�<��~|ߖH�Haxg�Fu���0�$��`+���Xa���o�N��p�8y�E���rt�,�)�Ė~�_�#uĠ�03E� �F��k�Υ�����	-�J��F$A�W�\��4�x$ �>=;ȹ��[�(2Y�U	{�J֋��6zF}�aT���.�o!��@\�5���ݨ��N�N0t��z?���7��C����B��?��X�)���R^��Ϫ�	C�.R�U2�B�ŝ`�+-��  &�ʧ#w�ŘO������Iv�l��g��'!�b�6@ᦁ<��_�J��Gd����c��`����N&`h�vdKb����p��������MEK=�̗��G�`��ic�������ί�>�x�(hp�a~���o�J�3w��e�����z."mg�!e���R+0�a;���I�f6�
�z^]���#���N��q����@4c��������o�x,l�Wq���t�y�N����"ؾ����L���!~ұ��G���.�@} �G$�;�p��V����]�>�m{3�ߒ�K��b�ʜ$o>#5�N0Ym\F[��w~��q"��O�+<I��%6%`.�GiB��ڰ�HZwG�j�9_���f$4�v���3��p¤����E �-�p�9 �c�8�_�"��e7ò�W�,��.s���������ݼ���̛��L�uQ��4@�I��d����r�0Z���Y���+��<�Y� ����g�@������ �"�h�������=�$��)0#CIo��`?���2��7��!�O�x!g��e"� ޣ��qČ�7�\{���gk���ٵ�r]��-��"��:�H��-���	C��6Xvi~���f�χ��޾�M%x���-��9BS,���d�V^61��9�b�~��m�󱞮
1����[%��W�L�sz�(��[�����6,����R���Re!�AM�UM�X�d�w;�bv!8��=�W߳9w�=B?pGj��X3��<�_ճ����Hv�pI�o*�H#�z��g�5_DM�:Q�'�j�6�X��J��W��ax�,����j�p�#��������� �VD�j��1���#� �*�6��4��I�?��M�S�~;����Z��`��)�6�(ej#U$�ĵJԨ��)�T@K��6���h%��v����l
���Z�� �L���A�	�L:���)��ّl���n񊇦U��m�r�TJW��d|�sh[y��TSK01T(��rf�Y�X��KR�ْ%����^BH�б�gX�Ŋ���nf������
;��2�LH�k]�����oH� O9g�
�zy~)�E�Dh�r���[GT.ș�����OvKqr	�lqsLv GQ��l���*�����B�
DA�F�]��^��f�YSӁuߙ���k^)��fm�:��/��+�V��A��֕�Zz%��X�b��cA��{��رo��N��H;汋8��-���8���*��	��2��� !�
n�g����c����8oP&�I\��!�,�����Z�9�b֊�o�%[��)&�]/�)[��ј����8Υ�l�D`4��+O~�ٴ��`�k�Uc�/�w-?����m`����6�]k�L_�0��.l���{ �����Z��H��k����~���u�7)���gc6�Ч���ń/��Nв�v��&�e����!t��o���_�����G:�f�8�	�`�ċ\� �?r?�A�������&99Y3'�%�VF'�8�X�j�fd���H�'U��m^IodV�觡��+{��<���;W88���:m<0X���P�'��O4��/���M=�n��״�i��&�Fo-6�����qs+�DO�B-6�怲|����~��[h��$��OQ�U�LƼ�� CD1O�o$?fR�>y��K"�v�ª���p�����	� �I,g���񁵭di9_:����U�GY��(��
���w~���ei�O`B���v��"U�>+$x���|���~�Ύ�Bx@in��g�״�%`�s��2X��|ڰ�m����3�s�a{���MH?��k��A�8M������wu����K��͟�j<V���4��<�ܟg{f�Bi��:��i27:9�&Q���L�kފ
Z���fq�Ŏ�?�As������?���;�ʾ�0��J�Yu��L��O���Ԉ�&7���3;o��<��4r	�$��%`*w�1�Q��=��c�pn�vE�Kr����2Ho}�v�!TO��,��.��	�̆�uح��1��X�������EٸR����@���������[=) �z]�{>���s���A�̸�X�"���2���e��(��X[�
��!�z�y��O�mȌ�m���R����6)���FV�E�J`��>��*��Kw�_���� -�DJU�9t"X�ɚRw�>����1���?�0e.�X��;�����.4��P��*χ�+V��yo�j>��m�� �FZ.
1NL�SRR!>���Q���{�!|�ϗ��\��
�?�[A������iB��'��'�W	���:��E�BV�`>����K��oZ�Z[ьv�Phe�$U˪�,4���p�?}CVG�D���Q��	5g�e#7:�w�o���6|M�I�X���g�O� ��MN��IA�zf a<�2hOK��=���t��H5����Ԭ����4`��zq�rvf��7�
!r�>3D/����S�9��IbJ
%��U��n'���ڶ��\
~{?H�0V�s��v6QE���Z�0�c\��F�Z��_-�;�y�v!pc?�Pˤ�ϥ�����Kb+��xbs�IaV$�в�z�n��k7�������G���t1{�-�_<l=N�.x�&�]P�o��+z��ǿ�{��:��A\�b �x�=nhx�n�Q�b�J]�ڄ�3J����<&*.1�Ĥo�۪V�tWI"��t;gJ��b�a�Y̬>-���Vl��|�����'篣D�Lc���ޣL%�<.�&�$MA1���	�������9��ȑ�ɇq��ڿ�E�"N2�߼#���F�حpR�=6�� 8�#g�IA}��Vy� ���G�{k(j�gL�}V��˰��[&�IJ���ۈ���|rXS0�h\����R�^g
��(��=��p�f�˧�n��{c������iZ�����\��:�����Ǣ�����}��.�������̼m�4t^�&?�)�����o�	5�;	}۪9�_.�C�Q�q�������%�{ �Y�= l�!�?�a��`�E�f�'܂{؊���,aF���aE�g��P�^�.P��BT���������#w�\����T ��j�qv��@ұN7Ɯ�:®���(*u+MY�؎G֊�c�V��l�6�=����]����64)�f�bx�ں�:oGa�����\��TD{4^#�B�>Q�3[�X�A�Q�=SKr�/o�U�ߚS��`�hR����P �=�R�"���A{�w��n�[eت�_y���jq���m�����㙙������7����q#ͺ��}���*�
�@�2��}�Z����ҹ"����ᷰ~��)��j��oA5�������ils��75"��$���I��W�Y$!1���-��m�*H�I^պ�70s���Wɐ�u�ؽa9`��/Es����>#� Qv��=�S��k�kG�_>���f_l�[�*z��P 4RA��WzM�ˡ 9��RK�=��i;�����������,���7Ӓ���OؠEx�m}���gK	Ɩ�l[/����ʆ�p�[J2���ߎ�.�FZ�5��wdt��[Lq��6A���42X�Z�Z$�yu��=7����'�/�
XM?\��䉵������g��3����;����E�LnQ4^�[� ���1r���a �Ҽ�7��簤%m����P_�j�Q���� �f��{�be_���,W9B��^�:���ໞZ##;�{D�_ �Q7Dt�<�Z��A��y���6o
�0�(�̨�a���Ee0.\�4�G�l�jC�?"Id�-�������ipxaƇn���e���g�s��Ң�W���ĵ��HU���d'BW]_�����g:*���������D���돜b@�ΎB���-���#p��{�[4�v呦o���SSqn���?����Է�����:���c�j)�@�Ħ�7�ҋ!=y����T���h�,�K3�����`�FPa�5c�\/��#���I7�G�َ�7�sL;�W�N��m�������u�!>6H��T�:1�&���.��>��y��PD�'�~�.s�~�\- Z}kR�w̒Vn�I2D�Bs�j�1&Q� tk�f���1ߤT�k�����+�,���W�1v�����������vbz����$�*M��޴��LΣAoYk���gl�W�>��&��l\.��T;�Bߕ�����<uI
����"��;�����E8|�@R�ld�(��*f_Khx�3�TRJl�"��=�[["60$����1��dO���#jd�=�w¤5�����"�knZd '>�Xԁ��d�N�f��>�Gf
0�>Y�Y�~Z7�7���s�3����`��9�"�Y��ĭ��\%/�l*��'���}lJ�� �<�0;��@5wOy�78J�������o{L4Wc���4u-/<��c\�7�����-��yS�Ğ� u�>��_z�}c<d���3��Aĉn�����g�|m�|��3+��γm�У`�Qw� �J�!E��򾮦��1�)�e[�����,�������f�[�l��Cu�R�a#��ڣ���^E��HK��; ��-k�̯�gK]ю�?���މ�p�kY0�5>��uI�K˧��!3<���-��؁�6z���/\h�w����s�	%03�خ:��e�~[P���O� ֐汽p��#�h�l��i�}�ge�z"S����Y�4���Q��Úfҁ�l�:����S��Y_��kvgp�ZDup�L4�?�|��;�(=�c�E��@ۖ�nG˅"�X�)���u�L�}ԻWڣ�ML�U�܍b�K�`��ڥᥪ;�9�O�`{؅�b����H�bAM�P���c�]�E���h#�'^\I�{�.��%�o�:��n�ȋP�9�8�Qh	)q����	w�Q��{V5�Vص���В��Y�2N>T���O/u|*\]��{W6�t�s!-���x�E�XGIy�L��\�e=2�I+��2���M$4�����o��X�TT�P'�Ji
>y���cgV�&(�M�;��_z���yi��(���XR{���i����o祝W�@&��|�����p����8�Bp�����,���I��ɂ#����N�It|:��naO����ù-kJnW"ݡ�O&�}��^J@2H��h��ɛ�G�>]��X<F3]ʲBw�����*����boa	��=1p������u�xϗe��ѻ���t�O�o����I_�� ��֑��J��:_�������rHx��	G���,*�U��nP��#J��2T��h`\	TUa�H��V�����ǤI)�J;���GSd��A�6�r*W��ɋ��VO��o�V��`��+��S��A�Vۏ��������"���i�Q�27��C��� ��l����ƻct�f-���r�+�u`l��,d`ފ��Z�6]�Ƥ����?�5���V�B�kN��'�ʰ���� ڪ}F�ߺ�\W���GĽ{�`�b<a�c�Q�͍��d+��\}�4�%���7;N����a�vP���HG���U/2x���m�O�G��c�5E�n�ǜ�?^�w�g��0�;F�9a��ï2�P�h�i�x'|M���)�#����a�+5:�q�����ܲge�|�gُ�� KB�Q0j�����f����}��4"�u�Y���z���/?���c%����r��.�P�?Y�2����x�?G�k�o}�Ј�cݞ���G�A5UV+c�r��hi�֩2m8�I�3�t� 骨8�G��<B�~G�,��=�����O�O��2�7�ള�A��M�@�W�m�2᫞3"�|�uW 9y��F�5���G)K*��~<���(��t/���;�i ��W�����n���ik��Xh�p"���U;2���pS�)���èp�Bj�UHq&�/Hf<,r��Uk�NW���!�'9U�ID�^���˞�4�-��
	G���Ҭ	Sa�b��۩��)��ډ{�(�!������E]y"U[��Vi���2~�r� }�2YX&
����[�6��:(��R���SW�����lJ��1z�5��MZ�/F�����b�e߇��ŵ�7/�����~��]Kx��}�#,��J*A�2�u�d,���H�`$,c�=F��TᣴT7E��	�&ކPrf�K�$/��u��{����ijK�vG��^�Y���؟�}�.��'o��K�+y�E�����Ye�x���ӑ��۳�]פ��}���Z�ý�K���O�#�v/cp� ��ywvӅ����JH
�`�W�����
���<ԙx+E���h�
�~�M������\S��Mi�0�ۏ�|����*��؍[TV��0�ԱTc@:]��J�E��[�k~i��q�؏٤�$�7������j{~hv�#iM����B8�_����un�1�Q'�(�
h�5���#�f�D���� @�|u��7�\r^��:Q��e�6�;T��!wq�b�V��K��Y_ �I.�d�� ��f���2m�8�#������#6�]�~�S����6�"K4��T:�[�J@Pi�n.��~�ػ��g�|DZS!�����̂����T�gW�5�w��ʀ���}�""�.I�z����;<!��2,n�,�n�ؚ%��i���@��Iy!����݊�2K� Η�ؖ��2|G�ꫛ��(M�DK'�w3X܅�]�םJPgOT� Hx3��$�\k��{��E,�����Gk<'\Lʾ_ރ��$'J�@O� ұ��� y�:S=
�$�L�1����oK�%S z�"h�[ ય�Zn��Ue*kpF�k���XU�����ܽO��3Vݮ�o�@`���r�'L*:��9L�4�^}�n��F:9���X辧0yޠ�� t!�����<Ǝ�h�y?�`�<�N;��(b�^	�
�!�=A0r�VƂ�����L�5�=b�a�ʮ��*��0`Ry��5�#$;���"��||�ʹ�f�7�!T����!4��P+!�/9�P\���e�Vݱ�B[V����*j�Lst8�
��ɼ�%"��K�$����e�DoW3���0V7C�Kg�a���4�(���]��.]�H�=�������K��d�.�B�����9�[�t��>��H�yX���9�!�l�۠�@�ڃG��8ȍ�\� j��g��=�����+��a�[)5���<ӭ�S���	2�aqzdS�N	(G�_yZ�\�T�5���A�G>%m���5���3�U��o{=[���ʟ�B\��ij�f
Ok�%�9 �D���ʌED�B}�~Vz6�ϗr�1T���W���K |H�n-[Q6Е��n�gAͳ\��0w�`Q��SYT�q�W$/Qw��5����$�r���P1���t���N ��;�V�v#�S����Ѽg'��K���@6�&ݾ1�oG�?����W�h��_bxO�聩Fu�=��p��q�_�sPYQ��;����zrJ�"��7�:����փI#֍d͹-!�bG1��r�U��Ω{�*y�-�}<���))���,�63�L��e4�Lkǿ��%�� ��M���%nd���P��0��?�\q��,e��r���\9�3}j���0q�z�
�ķ�'p���n�gS�ג,����S��c?A:r��Dg%��\������`�G#n;#��Z��\:|)���;�����8r���*`r��j���%�\�qPN�2�)�%���(xe�ࢴú1$��"�,�v-~'�����+z�(/A���[�99^���W��~z��<��g����
������3�i(y������Os7k;�rJ`ӫ�>�%7a�V�(�_)� xf�0�i!>nT%�=�S���bDͳ����b�"�?��%�ljf!�ģ�B�p���C�z�� m
�:|ɯ�u"�g�����58!�G�L*��f���ǡjǁK�W?�Kz]H~w�� -�k���&v�x�$���V\��Ъ�/��ٙ�g��`�Ό@q����玂��:�zB���g�oU������j��e��dZm\��k{{�l�}�L����S<E
�
i"h�%̆������7�VbBb� Rf0�1�K�~�x9v	E�>I�tK�N
�?5ƙ����_�/��*�rNS�1�J���OGF�:�G�A�rd�n���p=,fg���3"Ib��a������2�@ק�Ǯ P��`�nJv<��^AۂΒ_�M�ܨ6ս�0�.�`Z �C�U������CXgq��$��nɳ�|����m�-�ie�'BfQ�VCE\Y��3�1w;�{yzdh��Υs-[5)�=Q�<d��lּR��<� �㧠^�r���;"҂�Uj:N<FU��M��ޯ? �^Kx�c�~
S�m&���Q����),Fi����p����6vQ�w�2=ҜK����I����B:o��Y6r!ޤs@[�3����ߣS��Հ�;�e�!3�Npv���!�LU���!�\�ȉ/R�W���e���&�fE���kt���k>Z����J���e�.t�=����.�����AG׊��T��R21Js�.��U!��AC'�ӕ*�Y�P��y�lþ�����S;�,_��s�6RV2^��+�:���ƥx4��������l��!�(��������:kjI���c"�?���HId�]̷^�*8����8�MGQ�䗸{�i� �3�d���;Ʉ����ː���e��lg
�t�4]	r����b��-	Տ���CE��=�B�Izw�x@���?pR�6�%�Ԕ���*W��$�Ɯ���'����j�o��&n���#s`x=�-�'����|[jM\0�	޿��#/�!�b5�rG�u��ğ(�Ҿgc2�st{I-�6�i�%�bXm@G��\WO�p�ޓ�a@��G�N����s������Jr[f��u��T����g7*ڝE��v*�Gn4�bZ	 S�%��B[��K�!�г�8������S�X�֐I������KM�Mr̀/d���=�^mᘍ�I�I��7�ǁ��S�BN6b��F,�B��Z���ZJH����H`�լ�W餭^�S��b��6�T���ҋ%���隇֩F`����b�2�����i��#ti����mb*4��4�yܩRȽ��9Oc��+������c��S$��iYC�.;���&���T�a�R���]�,Z�j��VT����=�����ۦ�T�$��G~�+D��P�OY+l��p�5����C~����=������ߎ�nQ�3��6�����ūwd�8�\���o9�<���yejp|)�SM�����y�ߣ�u/��}G���j�2 �]GN
�yQ�pU-���q5E�f�����Z��6�N���q.�մ���*g��ui@M�{.��OV�El�B
�S��J�	��'�վ�H��� jOh�o^��۔�s����צ�����2��u$]�#��x[�,+����G��8��.K9�>���ZB�,��/�O٫�ն�/�����c��m���_�Il�f��쀏�'���{�ڴaN�Ľ����j�j·u��vt�Y5�@*fx~t�M�e����"?�^9�(��S�0VD˰V�_�u��.U�O<����z����B��u!�!����>��T�K�n䴝KF'm���5�9k�ߚS.of�^`�3�xl�������>��KS�TbZ��_Ӵ�G\Cph���@ :�������lc5A�0�;��uf��S���j�26�KI~u�e������C�6�J�j�n��w�[�����7¤�N<a�w�%����̦βjc��8�7Z��;5��,T*GA(�	��UW��m� �(ɩ0��6|dӰ3���]��4�����_��Q�s���<�� �G�c��-f�{G(-	�܋K�g����1E����=V�$�k��S/����=��K�_T�o�����,ls�n���QwEӵ	ٛ�2�z���w������޼�-*TC��O�fx��*���"�8c�G����\1�(E:��Z�.[��3�7d�;M+�U��5$T���stX�_��KN�M��b}n�٧}�$6>�@J?>Be}�#	WeȘ��:�����q�,B�YE\8�\���4��F�
'Ãɧ�`�P��L@��w�Qg$�SZ�[�*a3��4��q�yD@Fm��x�M�R�x~>����$
���j����M���|ݫ��y7q���]�jՐB�>%���
6DD?hM��3	�o[*1@/�8v�86�w���O���	[�)��>T&�H��_IEJ�<�B�Y��w���+\��M�K��
�A`��r�(:�!Z����%�>/��ER�E���f9ٜci�0y��q�� 6T���e]Z���*2s��i6��n�>�!f�F!�BI]����_P+�-�Swt��/j' Uy��a�.���R*��3��t.=��9�ے23��U�Q6�~!c��*T<GS�keU�����.;�q����]�a��$+ ��fI��n���K���wEa�9��2�.e/�#����g*�V���+�&Lo�ݿ~�NXYh�*S��Y����sq}[�[��|��`a-p��_m���iqS���ѣ�^�b��{@O#� 9�����0�\�)��%�o֪{)�|��Wr
�ư��(��h^fw~�{Mg)���+�21����(�֐�8� :F�xK���M�2���H1���Ae��D��ͮ�V ��B3}4�F��;����|f�a	��"-����PyX����~���D�q�L�s=�G}�l�(J!y@{^T�X�v}�9��֩)T�2�J먨���'�{�4�=Y6��n~�@�&���y��I�Ȫ$�#�7�-g�����4K$�\6�"M�p����G�M+��hK�ܘɦq(�-q����3�	Ä�|�<ħSֆ#��CL�tK�y���8�>�;�mv������dh�g�����[�������� ^�~O�te`��c���<�wL{�X�8���8�H�@�G�a�LW�\gx�����ͯ��i疼�P�5�O����j��;B�۱h��>j�C-"����I�^<�S�,(�N��x>)��0��h �ȬD�{G�׀�~f}Rˎ�;Ӎ6Q1��_ �MM��X�m��r��b���z�j�ԹYp�e��Dznbn=;�E�#B�N�-��S��C��N�5�|����$��7uP_�̯=����T�[����ǜZԹ��w��ĜY��~����>��fRasu��V�P�C�h��6J��6�������HܒX꫻�P���V�J��O�m?+���\��ɍ���$��G���=7=��0�=�-;v��7��:��w��H�ԓ2˟������I��e�OHΪz>77S@[Y���� ���-��-�+��ģ�Vͅ���1g�͚fZ�L���Ƅ�Nگ�O�w�¿8�g���w {\6P��b�������l��6��W��w��<��R��L98�>�R
�9���{��koOL*SX���Q:W����9�^��!��:Pq�ȢZ\��qC4��_�c��]�ȥ"DBl��q�ق�4q���������P��Ahu`�W���
���6���M����2#N���� �ck辍�r�̑��t�����>u�F�}n�EѦR5�e�	Qun'�S�t<�9F,���$ع��v�{������Y�?�2ڃ-�3��Δ�gJ���������$�K�tn�@�]	iG5r7E |˥�Ўeά��&ê�I��[�U��S�x¡��i��R7����-�ŭ{s��2��WM��Lh�Yo�9fG�� ��?���%��)}i`PH�*U��o.c���^).|��C��@��kTA���M�HR��ꏩV���%��9� o�t��ZDR����~��sx��Ct����GT���3�(��|�����G?�C�|kߐ�R��?��f�/we/���x���>�U�w�+�Ȱ�������+����b��>[�z���J�gp���B.f	�,�g�Ѭ%JǊ����1�%��6˸1G���zZld*�h���*	</�l�/L����C	f)��Pg�E��'[��a��`KG=��0aZ��3ⓑi�����T���\B'q/>�WMz�ۅ������:��XL��M��8EЮ��/p8���7�y��K�F�u6��J�FL�=%/ٳV XV&�Xn.1���8W�� +[��U�:cQ�U1���TXtr� �HB��>�֦�ُ]kk���VG���E&v��@ �����׸Q\��3� �2^-	��K:�y� �>E�̱��ר��A����ֺ��/�t�
�J�� � �71i������U�� ���6�s�>cQ볽�����C�򬈫P��5���)ڶCDnf������ƜO�EP�
A��3�����������ڗ$���@Fy�R�&& ���+GR��x���#2 �����ҍ�0[	����k�Q�5�,��J�;[L�����K�>��`-'�g�-@c�u���A|̶*� �ހ�B�=���z�g�3����\F��#����%�]�'��Ya�Qn`ve�����3+_���G���y�!�7�VĻS�LD�S�	z��4�=�:M�m� ��AD��Rl�PPl6�����VF��:�$�ǡ4�S)H�;fxE��+�����V�q`M
�U��ߙ��@�8�>|.�z�k~6$p~�
�����{9�)�~����వ���< 5��Vs��O{ax�?k�,@+�����`Qn'#?+(P/DK�jH�縶1��f��o�G�W$/)����T������%T��E/�.g���Q���@��.Ֆ�PU��N�W���Kﺡv� U��먅_��6&�"T+}Gܩ�WY���t�����O!���%��3,��~��X��t�m٣�4�7-����:������խ�]
�GuA2V�.�v�O��A�ͬ:��,����V��u*}�}2��!� �/�N^��m�ç`�=�vZY��gV�!����VK��*�/U�sّ�qt��&g^C��9`�X6�����U<��pl��083Q]��.�6A��8 ^J�f��0�m�vA�^�����r�.(�i+�X���B���ɣC.�>�u8?����}.�rH�]­ՙ���J��Z<�
 �`�0P��?��X��;g[�������u�lԩ�5~Qv��c�*�_T���{Љ	��c�E�Mpou#��C������Es�?�e�-��b������Y��3�a�K�o�얒�{Όa-� �����ِ&�2ZnA�9ݿ���������k��0��4�Xh��:A��
>��b�v��M��DɈ�F�W$Q%�&s�.�p�\�9��Us[{��� 7K��Mx�_�L�}DX�;�l�<s�c��f$�~x�uxa
�uմ�ۀ��`��S����)`����{���$IƬ]��G(��Ы�7�FNIS����@&�Wpb���+�ɲ��o(�'&p&q�3rA�9rV��buR�d֭6(�p�3y�8�s'���
sF��b֧-wb�_lq`��ݔA�ғ@��'d��n��ǰ,�����t�t�ȓ¬۵���AKQ1��A174U�f؞6�gfL�w�V�H��l�ȶ�}�T��a<�����F �Az���4�u!���<R��k�ᬛڝ����?N��H<�P�c)�8�XH�p��y���L{���Ó�a�#J�QF&�"UF������nW������ݨe~ή�d����S���T�V�cP:���r���z�%�[�RniZ31�����jb�پ����H������,(L�"1�(<�����'B%�7v"�`�~����[��*��I��Ҙa*��w�R�O�R��c��B�Ec
*�ʃ_�(\d���Q���>[4��� �O���ȉ�yc[��lozn@���Ggɑ7D��%�2��|
�aJ�W��k�����`�I�s�V��K���a��L~^�#u8#6W	�:����w�ewKF���o�F�٭1��(��_m뺡\L�x}w�sG����*t�R��
D�w��a&9��),��M����X�B��`3L}:�Rk�U]��;�1���f�vu&Ys%��e�j�=�3�����υ�����[�JO������5:��A�',�G�^�p����RZ��᭨@p�RS��h<|�?[w���wmc�s*ϳ�FB�d��������N\��3]��LyeP�&]�=ݜ&�f��Tv������{�-�g�'��Hi㽇�R,�[�V���sb�����\l՞{�-9�GUD����T�z�`��>1g0�~���qW�T��ɿ�pmÑD��$��4�v��#՘(RU3�w�[6`�ᝅOG�i&BW�Q.h�8aX~7^�=�U%[(��ѐ�Go���4rj�-�2�)M�K�⭩&��L]vu�YGs�m�j ��Y6S�|C�~�=�\F���?�����Sl�!b���]�Λ^���#�<��]^:\j��s�I�t��'�6���Ǘ�3'ָ2��i�8��x������G"t�^��
 ���_��	�s��[����Ni��b�������5�f�#U
�xs!;�
2'e�է�F����R���������=�Cھ^�6��rd�\�P棦��jj���1�Б?�G�o
8��p�=^����% ��k�׌ޙ+���J��g/�Ւ�q�a��x,v���� �{QC${�<R��.��gY�%<����*2���je�0Ě#�P�mĔZ�bTZ��9p��e�O[�ܿ� �i"\EB6=_���2N�p�T�e�?稩��3�ڕi^=	M�sED�ܤ����I��ea��j���^H����*ӕ�z�N��(��{�\���)@&Uc��H���xk�
ȍ�f�'�+9&&��M�_I�K�y*����/Ǘ� �jj�������/������KZL&��e��)�L���2�)��\V4u$N�s�@��	=)��C��T�HDQ�1ݮ��f5ˀKpi٭�tN�?���f@�n�K�ٔ��5�|%���cS�&u�_E;����ģ���E��W���Ą*mC]�;�z�<��lO������iK�SBW�
�ѵ1S�&a`��8���syd�$�m���`>��B�Bj6�F�X�)���4�Q���'Ft�6:nK'?��Z��_Ƕu�d�6q�<Q��k�O�_'M���-�)�!�@�al��` .*w�Vڼ|�޶Zu:��C���e�9�V��z����䖌�f�t}�Jt��؇^�����;0�o��ơ������[hp����3H4%l���T7����~K�xڣ���隻���I�P�+%+��#����;?՚tp����L������L#�քbʤ[��bc�a�)��`�ƍv�)
xL���$��3���ŧ�K3��}/t����W�7���Gk����4�.���w<oG�}�/'��Ԕۭ�D8�o"���KCA�>�E��iUkM��V}+�8�dH۪�>S�;�ȗ��../�S�@��O�E�����aB��2T��n��?0Q6���
�L�F=�>�X�hp�0g�_[�%�&�j@Jd��^�j5S�o��`��X��NM	�}ߗ�����q<��P���ҟA�:���i�J��+�����8���=���,�D老mQ�|M\��,F���|�o��:��3���B�N'��|�RS�ѺO3��,7�}�0	Sh�>�=��	'ŭ%�ZP����JZ���!�bg��(�È�rta�7���80%�f -���#�lɎ?��3~SN�`���x��1��nSNG�;I���d���%�;�mq�v�J�Wh�6��yA:��Ŕ�N�\���8�e���}а��ϷM����"�k���b\).�e�8����� jڤ�)J"�d�Cb�$�c"�=ޔ�+nՖChn�i�e�V����%}ȅ`��K����~����e�XD��4e��B,��~�E��:�к��̮�\�h�P��٢��L�DO� ��N��c�S׸�!�T�'��6�=ֵ��(@Q�Q����az�eB��6F,���z���#-`LX�Z��aR���3���?݅1ſc��&�{��\����>�4��Z;�P6��e
�2d��>v[ ���6,?������hK�F��-��_���u�^A�J��/�������`�	�U��?l%���MxVN�F3
} ���_Y�M����l��نʾ?�W3�+�=��"�!�G�")�}q����:��p|�*�|�s����ٓ��3P��0�C+���\[�\����/�sb`m���)spDF�4^���kp�?ղȜ�k��>�ڴk�ƶ���^�}�.���n�-N>E5Y��|M�c���Q���&�ܨ�bۡ���/���`d��]����e�u���|Ip.�����0��+a{Rpp��8��'���6���W�Ӈy�#�����i`L�^��%���d��@:�4T�0�u��P�~r��frO"�F�8� ���4�Ba�*����F�ݥ$��f7)���:��m���59X̌�i�*���#T%\ӕ o$ή��7��a�R(�pNW�����ru�U�꿊7��ot���m�����EF�8R(��Y
c��u�:\��B=�����R��vB��k���UV��`(��,Dno!dO{r��"���i"81˟pW\����`�Q�賈`������}[��Ӱ�E%A��4gPK��n���β^s�-���V\�%6T읎>��X@�MF�O0���Y�r�|����70�l�SQ�Nn�w�@�zū�[lG��o��<�°2�������"����[�ւw��	%˧��)�����p-�n�ŵ����4�u#hrQ��km4�����aTsۥKq`�8�Z@/KK��GUҽ��s��]���O�n�t84)�Br��s���D�C���\���ֆ�ZNM�r�_�1]��׻���l?���[n���~�j��u$F����d���auL��Z���Ġ� I2��_(�z��3k��q.��	��gޠn��H���+�B[0�J���%�T|u|�p��M�Z	"���Q5�?�o�+�\z��P�%;>�w,(/P��<�=�������v�8-�k�RAh"���@%��󎤬�m�)��j:����7�/���c��F:/���U:3X�^t}-��Ҵ GA�����_���e�"�>���+`��;g�X��ޓmζf7Y�N�!�"^��&Z�����ٿB�@w�M��T�*�#���h�C�<��� ,�Nˠ��k9j;hi[T�V�m�aZȘרCl�?�hx����JFTG
�(ԥy=8X��+�����شJ����58,I
���/l��q긓�i�mf�B�^�Y�cqq��F�ED�7��="b��q���/�X�J;����-;<驓���������5���S���6�+/� �'	*+!Yy���;��9�qd��#������SO��Ї�w"�:��n����)�1%����|���;��S�h��CWf�`� �� �)��$}���&��=�L	�!{P ƽ=T�� ��>�o�W�&���������3�� Mb�f P�/,�tͤo�a�<o��;%Q�Y�46�T���6�Hi�r�N�>K.�L��h=�9�Q�V-D�&:������1O"���ypx��Mq
�Eb;r%��k�I�;�V	�u��,�ALۣ��<��?��]�9^Q2�D)����'31Ň�GL�.�~Y���K��V�,��@��:H%V�����8�d��e)�֩��e̛�t��?�3Jh4{���'�fsC��4i4>�����u�ט��_m���_�0Ee�2�s���<Bemw�PI��$�*���%�fZ�Q^s���GÅ�٤c�O�~�w(�I
3g�}��Z�e��P�˳⟏[�t��/�,]�/��I��s�l"��� �]%��F<چ�d`�.�N�EHԉ������HdG[���y����R�����\�|FPM��K'M`��O:�"b$;8��T�IK�3=����t���~�
�&�����V޿IA�hZT�Ƨ;[ �+pf�&`Gc�4@m.�w֗aS&PXV|�2� A�A20��%�d�j&"����׫OK��� ѳ4HIte��ˌnE`]��m���x�
��Yp��S�&�aUbt)��?�u���& �����xcMT�i�����L�稱�0Q奍� �S�	��pj7��x2���in�0M���3�l�����hA6]t�M�y�	;I:�5�/���Vcu4�Ϫ�g_��F�5Hy������p��Lӂ�Zk�8CU���r�Ui�r���p�2.��\wp�]��y>G4�q�>����"�����d �t��FV��<þn�HL�-���� �h�3Q7<�FN�KY��'�f���%�a.�0s�ҧ2�|>����3��;�A
�[�a���m*h���p��ɵ��[��R��������������3��C���o�eN3�+%_��b����V��ȉݯFH��.�w���d��I4W&��/��� x�!b�X�����$�짝��x�k�G��W˙�]��I4��n��Hj�%
�����F6��M�J7��{�8�k���?jNq���@M�.��[Nu�V��M��ع�I��.A��\v
B��n�E���P���ϥ̥����.o��ҷOx�hfl<�G�Q[����*m�ܳjG.��Cp�*�Z[$����-��L��`�|�Ѝ������KFy
��}����WC�$�5XX4Լ9��>�A�5������S��;c$���!y��fg��{���e5A.ڈ�� ����1']�9 L`"M`��F��괙�x���Fmt�Ok�����������9�0,qL�H�L��	a��@	�J�ʯc���xKn�p��)AltA�8�E�A��RKx�$^x��k�	I|� ���`/H���usQo ��ř��s��öy�K<��"��b�D���3�qf�u�*MG;o�A���`(!ص��+����[03MR����2�=���-$�C���E*�n,9�;>���m\��^5��"t���.�{V����T�ǻ���]&#���=r��Q�O�倳 n6���yJ���nz����&v*Q��m*�z�ۤ��UY"K�kGi�q���yY�W-�ӱ�Sm�y�ߨ,
�Y��Î&F�H�`�_@y��:Xcng�O��.�o�P���GEQ䓣��O+M����z�$�[V��ʃɇ{�a{�Tw�>`X�7�ʑ/����m6�Δu�:���`�y"ë�ٵh�4⩾?}� ]���AbW�X�C��6���_�aB��?	S]�~�ֈ�D��Ѐ�	� |r�:^��jя���(���lԗx���Ԛ�0�V[~�|��M�-�94���`RLq:�`M�h=�C���O��W������ɩ�FJ��VfY6[���T �J��TB���1��B����)�ב���\tr�!�{-��,�Y���DX쳹�Gu9<� ��v�?��p��Rsܫ��R�>ςh%QtPDX�	pK��]�J�/�� ���/ǒ��.���Jz4�	ђ�C�0�ƀ$�z���8j�+; 9�/���p�.�#�x�UN��o�'��2�>�"��D�����#����g��(aL���Ʋº�k��')�}t0�k�6�R����9�q���Uqh�Y�R���pֻ3Yy��B�h�
�Ru�l��KG ڴ���E��͙�3�\�_䷾*�V�gw�͌�z�S��&����ggw%q���;�	y��3(w�c��_'u<�{P�<��L����;��gs�̈�)�W՟�j��'�Qm��}�9�����q"�:Z@$�����2�&�J5�n!��V1ggݗ���*��2�
OS7^��2������q�º�G��^���ȗ��P�dS��4vSM�E���q��&a��s@m8��u�)�E�W����wؗH*fAȚ�>U�1�n��	�v����<#A��2Λ��t��Q�7n����F&��p�ӐX#�
��Z��Ec����5fB`[��݉��uc1�#y�ҳ�}`>zb	��{#�*X(�	�\x? w?WX~e������P�|���u��o^��U_�hD���d햇��VJ��D�=�vh�Gy���>�3,��,�~b�%\P�ƌ����R/X]��L-7z�<;��P%J�c����+�	K�-�0�1��
�m2<h��������
�⸘��F�4�� y�Q�^�,y<5�x�{aJ��[1ɥ�l�Ӏ[�s� ~���i�,v�Xw�D��Ń^�o9�m'J�ư:���I�f"�����^�4k��T$a���u�qґ�[3'�WOx�x�_�|�T�I���$2^��c���G{/��2ݣ�7uR��OJ���P/��=��'��<0'n�ٖ�?,xە�Lx����{���=7)r��;�
9 ������M)��m>��j�]�@��&�^�@�����ER`�"S �����u_����_���ۑ%y�a��D���%M1_@!��h���M�1I��������H�����(!���NfS�!��Z�D~�P�M,��u�����BQ�W����mӶn�x4��Xb�}k�w�V"��u0<5�H��`J���id�-�:?�H�}HJ�����%i�G:&���N�8o+�����GB�q��<���]E�CO]�}�-���|3WʴC6��L=v��L�xT���E�����7^��y�NWg:��D�A�>�d�`uG0��8)������ rG�[��I5��c�ޥU4�
O6�;ab_�J�X�l��%}<�m.��ծѲԥ���k6ޭ�V�Հ�Ф����S1+��Q��r�D��t����$'��<��2wd�ZLb��}�5�����*��,���k[��.��#R'H��RH&���Q���U���/"G����`H�ňw���WJ� ��U���d`L˂� �b���$����Qނ�'��^�k��|.���8�A:9ܫ�]�=v�u��=����@�~�����I(���1}��ѦrXN~>р-�OBd�u����:����S�d`�W��Q��.���5����n�>�ӧ1u6\Ap���Y��e�C�`�R����ґb��s����ı���K|�v�TP����"S�=�!��o��Σ�%!��n��j	��B���_�}�S"�A��������?��Oj��/o��$<��{|!	Q�=��h�Ⱦ?���p�g����jG-�iQ����s��
&
d�D�:�
���,�Y�?ǲ:X�, ק��֢��M��s>a
�\���R�2#'6���M/l��⻼DTQf��|��%��/I��!�4V�Ў̣�.'�� �l���saW�ҿ�[�TM\9D�Ι���4)v8T�Po� T;�V���U���{0�ZT�����;��IIl���������^��P'Y���@R����.�����������:;=Uq���UB��D>ܴ ��01�3�t &���7��]c���zS�>AF� ��#4$Bܴ�Ɋ��(��V[�$��J��b�M�G	�M�τ��ZM�[2���ǖ9�G��q���g��!�sa��ٯp������㩪Zܭ�
��)��庩9�[X��;G�̟jQ�9�*�������+l1�!� ��\p&dj-�3��8�����"�ܧ�������~��MJ�8N@���#夔�濆�����oe
��2��@��L��E��r��w���?��N�5S��h�I4�t=PUߩ/
Io�Yj�V?:�Uz�4��ib�ox�g#߃��� �\�t�4M1{I �L�,�0 ��� yKb��
�@3�����������?Kֲ^kh���m��:�.��L��ҬkbM��Ǎ�A��v����t��%�8���"Ȼ|��d_3����?�L�����%��vyu������~�
�6&ٱ����^4���Y(��-i�e3���L5r��������VF�ıjG��kT���K���~���)?�ljn�����x!��\v�/#0wg���X�"��Xd���$)�����~ē�*�0��yP�q��raR�9�� �155�R_�Sl\��jhr�ю�o	���]M+I�f��Q^ƽf2�����*7m�`w]�WpK(��c�jOQ��9��z��nI3A���[���:^���B��
E�ٸ6�[��*�{kS5�h���n��A��f ���Qa)��5��w�v_au��5��w����&�N�2nPAu�;���};��$��ﲆ-W����Cb8�7�S��&�>m�����|QS^������d>���DV�=5��O%�u2�v>��^�I�6t�7�,�?(N�BJ�m���dW[��e���سK�E���3��~��!L>SQ�1���?���ƕjS˨e�o-�6�~�u�xz"���g�k�~luW���IIW�`Ű}f�18� Z:L16���-\��-�����x��T�	&��)�8Ɲl���*�?+�8��}�=�#�D�!ӱz���O���N_<?������_�}�*�I�Dڷs�}�^2`�����
�$ ���&Ln��
{�E�ݯK�p�ǡ�XȉC�Q��Iu<�x��I�6�pT�vA�Y��Ce�,�l���:�/?6#Ut@�����}��� ��Q7 ��޴yg��3�+R=�H�û���%=/�,L/RTd��PM#�k��$\���S�=����}�+�ݩ�	��Y�V[�Q�,���u���Tix���w֋^��w`Xq]Cͥ�9������5<�{q����6�=P�����Ӹ�8��6��,g�Db"W�3�3:��+_7ę��=���~X;�k��v7�A|'�������H��!�P]�F�.^��--r�2^��ᫎ*�Bm`�@��N!�a��h�&���KXRA�r��?K:+�zs�i��v�rtՕL�JPX�ͤ`�B�q��s��D���$͟;��$�����hr�3ZQ� {W��5_ʓ�O��fɴ��2Ӊ�2tUS��)���,�.b�0��~�|���J��Z���w�H1���M���%�y�:S��6�a���a�]�WG2)�L��,w�	�!�=��V���h��[`_�pb ��j���*�!��s���[G��|X�H3~)���} �tM*�!��L8�`��ˈ!ywGֽ��S|<���tOB�����ΓX��/}�2��"���B���4E}�y�[B�B�!؎���\ўI⣒d� $� �_�ʳ��[٠?ڿ������)x��&+���	�@��46���Un��kjǤbo<ɉ�A.�oA���)��@��ԸP�W&c�W�ظ#���\!@w�"TL ?�N��&A��2��i��a _<�S�`��<'�;��h,b��)Z����G~:s��6�����8:�K3�!��(��>,���f���0���a�i	6V�b;֫���I�������{Q\�U�( ������w���R��f�q1ߝj�K��Z�0|F�]��]�J�Cl�:h���|���Me�5W�~t�I�:1��1t~�ᮤP|�)ȳFǭ��.{�@P0ryxF�W��"+=~� ����}�4�{Y����u��5e=Y�x�4�����.J���Y��ŏ &���h�^އ@H�G%5z����(Ӑ�7.j=<����?K��Jo<K�^��eAI~������&`��ʬ*Į���;Wb����	3A��JN�J�5��T Qm�-CJl95 V>7Y���_۳�&����|�{jm�N��a�"����;.��}f�1,Z��B	��%�AD[��K�R5uh^�J���]z��(��R�u�+ 0�	7K3Q:y�GI������2wNxIlSj�������Uf /M���:��W�)Z�X��Q�*P��v�}��-�E�F�f$%�*��p�>G+%��ޖ�\^�ׅ�vDsl%��RNg������������=�*'�ʠ��V�GV���N�	N�^͉�Cj������l����({�3
ɑ9���ڑLK+?W��|z>�̧=���cf�K~���f�O-�o��f�5q�7[-!�V)�r���Q��὘R�9
l�|�^�)Q��t��&�V*o;��V�I]�e� H`6���[��z�߭�����+R�t�ƣQ���r���8��GÈ'�M���>�;?S�G!؈�`�y��YI��2ӓ{�T<�*��:K@)���˙-}��A�7t�qR��R�NIҢđ$�n����e�B`�����ʾ�-mȔw�}N�M��6[�8 �=ywN�FLv^�>�oeT����cN��.2]D���F���� ��6��Nd8�a��*�����{Ȏ��	|� �{x;�\�u	���h�S�&�bL��XJ�G⊝���(�۾��Y���
ϩ�$Wn�'6�< ����e���40ش��;���_��)���GP���/	a3����c�sf�+n��ʍ TE��A]��X��x.>�Z+Я��V!�sr}��3>�2m����O��l��ε�e�����c"�^1�Ĝ4�#�C�ICV�dC�=�3iًʕ<c��)���,	=�;�5 ��anI�T�C����a��>Wq��"��`��E�G��m`cND���/�G���l�eݜ�c�OoO���Oy�.��	���]o
�lh�D�J>v]6�XJ�)���;��D� ��`�faz��j=�%j]b|M�/Z@�W��D==T:E6-����r,E�t���Wm�Å��{���[PG(��O��p�����7 ���=-XI*]�<���3N)�as�l��7����cM�Mj�zz,	��f驏�0rh5xF�C�f�L�zc��n��B'�֜���}��s�
����Lx1�0�j�j�?�ouU .鿱/�A�C]2}�i̳�`�yQk�enA&̿Y� �0F}'n�$�у�M��1Ͷ��Ƅ�В��	��y��ݠ�C�4O2���v�QJ���&5�������\m]ן��
7�Z����/؊��X�Bؽ��r^�ԑ �N~m֎��"�Hƥ{cdb( 8E�IΘgc�謶�f���*%J��2�x##�>zF��e$����v�|�.�;g�;��(��S��2��u5��[]�1��1Y+�E�R��y]P.��E	�l��7!T<ȷ��i���j�<*w�w�v;����;�a�j�Pw�2YD��^x�_ˮ����&SZ����q���|l�	4N�n7�5��}�I����D[3dy�B��d�i����4�_��ٌgVo�������A�"p����/3���W&�](~:m��sK�!���� *�X&/S����G�#�����ӹ�z���!��-��z��Q�9��#�t��.MA����Њ���������]� P#�7uu� 7�;Þi���@��+�2BT�L�_x�t7�٘�t����?���_e�o��dD�����b`ktb��C����'I��)`��E>J���T�fT�Ĝ8}�����	���];�������U��`�l;�]�y��	pEZj�CRE��6�U�����ڝ������� ��52p���Ɓ;��,et�I��>0T�N�4_��s�a �"m�5e�E�}��=��{l�bpy[��6��X��Vǆ�JU`�j���\�y�$�"djg&6q;��έ}\������烜d $�xV��D�~��U�'� �wXW�����2�0�Ol�o����L�Nl=߬�@Z�!���t�'R��Q��'dԙ�Is !UZ/�,�����b���c��FX:E*ݯf�a�\�'��GG� |������S��ߦ�oB���!�4̥���
{@ss���p�b�\u�C㈀���� \���Y��h ����#���}�����@�h�P� V"�9��m6�0�V�<wp����*��sJ��6�O���
-���@p��@��U��ߎe���uul���^��͖�QM�	//n=�5ֿ��$�N&�C��Nc?C���)�jׂ،~��g�q��v��X�# qH�r ��u�	WhC�t9�j���s��C)�J�a%�byF��-�wZ_x���K��o�Xs1��:��x�RO�u�W^Q��XY�7�m묖G�;�yޟ(�߬�P�a�)#j������\����5������_���M�,���D���m���,�Eq�������}�#[�2/�hl�(_��=zX�"	�okU���Ѽ�Db�Y24�Y�ܡ�D<L^*o���S����J>'zd�ek��&�I�2�Ԍ˴�?�r���a�ipzyDi���+��qMwt�k��Z�OvS,��'���:��C\���Y�c�d�S0���xx��f�B%ƞ� �ɟ�!%)�+��h�$�P���X��]���+��-yq}����=���1a�%�׀�+1s6uފ"�$�oD���OK������q�t�=���mr��N?�����ֶ�n->��_+�B�����C�q�y�c P��A�>�M���a͏������k���$�\���/pr�&|`�����`H�q�x�|�})�k�`qUFt�k�^��I��Ɠ�[oٛ�n���R��ԫ���w3�ʣGݙ�*/u�&xm�Og����(K�p��ͫ��*�͐@4�bE�>nWQ��k�iЩ����L�3�i��Z?���a�.�{c�:;n�f��O�{T���d]��EG�=�X�@���BoH ~���h��x����h}���d������M��C���_ג�N_�c�0�{�?��O6��βɮWK���	<�����j�ׂ�-�U��@-0C�K��O��i'\Rkm��������i;���3����J������o���� ~�Y7|�ff`������P=û�῍�L6oG7�7J�Q.17{�K��E�8��������n����|󖢌6A�$�w��u��W	n�v�7��Z���%;�������#Z�:2��ѣ�-[���f~"��n�Tޗ�cV�)ֶ��P/_�N ���h@\����y�ykkt6(ۣ5�۶�:�:�MѮD[�_�,x��M���<�"�&�O��w��~?�k^&��<�S�+�0&�=M��ߢ-��c�7�y�n�k�)� ED���N5�Qy����t�2#�S� bs��Pe�����Vn5�55�ͥ�{m��ʦ�VY��5/��|�S��9�`�$|��/�m�Q�T��a��Z��U�k%�t7P3�y|wxr+���5��pc���B��	���		��vː��]�t36�@ЂN:���!콦	U�|�r����E�!��wn~��S8ͨ���FJ�$�Cޟ[Y�]1v?\P��#oo�S��)��?x\J�'�$�z$e��}|h�F�f<�4<Lƌh��J/�HK{EU2\�j+2�u7Deb�B�Ojk�=��Y��˱c����?�*��D2�URA9q���j�9O�b�Ow�L��W�`��f�Y+`�p�l��a%i��ƿ��q��i�f�ٲ��#u?��$B~O��WD�\-��V�,%<)N��5F�9�)��)��h�I������D@�q�p���Y�Ka�K�輇vO�ք�B-�B���qx�`#�
���� 8�~���W�W�	��k� ���e�_Ɋ�m[���,� ����K|�E+;���q �.;keE�i�ᒇ�
Cό:Z7�##>Os,e��X��sWyXW�?����+6㆐y�� Z���\7�x򒱠��u�m
�i�@�`售C��<�Dpa�Z����P9�i{�֭����Ý�9{4)��S�`)kޔ�c엿����:��k��<~-��jڼ�,�Q�-h_Q+&��m�q`��k��џ��Wd�W��Z	f�O�m����KꨎY��Y�]��FIq&z�����\0�(�2�R��mM�Q�1����ďm>=�D=~h���R���}�0UF�_:a*�ݟM�1��c
F[����9��C<��C��[e���4I��UՆ4K�WϥS���69�|���R2���.T fA!�Q9�2e�Q#18U>�D�J�<�O+Z������1Q�:��@d "9�uN�r~�
_z��Jċw�Z]�VcQ�.�`�Vqz_M�}Ym�owBy��fC�ڎ"	�	d�^ڨ��S!�L���ǰUD�p'UA`��w�
u��]��eǞ�kxQ]������n���.�a���b��z0�����q_��[@�r0��-ԙf#���ϭ�P+��9�2�v-���aw=���������_v�lo��;��Pl���{ ?�$�Ȉ�ώc��CZ^Pv+oA��% ��p�
A�Ul�8Hý#2w�qI�0���恵G$��{~��O9D�j$�lH���)�X�����-H\�
T���P����걦Aa���!�u��B�B����,�%uq�H~���a��i������fI0���)'����r5���Hq�߻���ݭxې��p��Zq*�m�/���U��QBxve��G�)�J�SXҟ�DeK[���D�k	"���,cv��y)_]vrfI/�H,�VR�t����,8�Y1�E!����eR���Xh���4\M+0�k3ݿ:6>�k#A5תUQ��$ ǲ��z��}��z��bW����*��/�h^�� ��A�x����-���]�P�}ݜ�S&f�Z����ad��e���i���|�Z�u�����[�R&;.��>��-�M��L"S����� _Մ#�2b�|�R߼�z$�'D�<["�P�N]#k]��ֈ6Fz��=w�q�i��?@ ����CI���������E�'Z@�e��6��Tnm�#�[a�&�)���`[��Õ�5Ys�ٺ';Qv��nym�� ����L��&���n�Gѱ����@[�R���2���x�sG75�,��a�\�s��\Z���@�&���^��t�cۅ.���"�ا��;A΂/���ބp��L����b@4��ϰҞD]mUU��9�ց��������e�[m�a���ݵ��HJ�2�F4��S�\j��̸�f��a��	���*f��|߃R���؏�B0
����~V��T���&�na����6'��GE �Z��g���gI�v8�F�ɾ�Yç���a�E��p(���Hr))����r]M�4�E%�D66�.��呶�G1��tq�x���Fq��[����4T&�~���/sy�^᷎qu�-���<33��yTĦ�4{�p=Il�֏C�z���r�}�K�@��C���x�������q|�\�ƕ���b�vK�(���CU������j�,��ck����S�0M�����Vv3bz'Kd��K�G��F�-���i��� Ǹ�ץ���l���Hz�<Q�Sw�����9�7R[n��1��hW��WZ�E������r v��!z�`(
���r�䜋�9���,Q�^�G��w�v�؟l���V��*|��@ �VQ����L �-!��i:7(�U�c�qcC%S�r%.Y��y��+�5w_jZ"h�f7C�+_�j�<���8k�O�h}�� �>�Re=6Yr˿}�fM�ۛo���B�Y���l^����N�����$Y9Յ�.S_3��<�ܜ�L�����M��d�[�H��1�4(��&8F�qZ���ޛ�f�C0j��D�d�.8����x�Su89����,�h�FN~�cY�� ��hr��	�2�ȱ4]_������W��Zr#O��-����`�MrC� ��n?8��%���@�.����8܎2��?^|�}xw�E������a-{�ʃ��lQu�P@i48=i�M��i3�1W��p2Q3-^���ᕿ���ei����P���B�����<��2w4u}Z�Y�ǃ��߀�{
k��r��.������CT=�X��e��J�����ثro´��������3
�Ro4�2f8N~�d�Z[ OB�#H���[<W����'� k*�����x�t�t�{u�njW�C�N�!g��n�uD��-�n�sձ
g�����ֶ�����	A~�P�+4����n�J��@%��Ij����qa�m{H�_�/cgk�GZdIN��| g�#��Z��l�ֺ$��� ��6%4�����	7��b$��-G	��c�FJ� SLTY�~3:cӌ��Yڍ�
��E�{�dʯ�m�~TAhHz��H��:����ɶQ������=��c�A�}�C�]JnŹQ�͚���*t��'��Չ_r�Ȋ>+L�m5���b�+,�g�/�,|�ds"jr���֎P��㞫GS���\�%-ס�p��還�o�����)�w�˃�:ӝ��iϕe�u;��)<�1�"Y���R �*ͬ�e�ï ��q��o�{��M�>Y�JP�	w���]H�.��c�%��t �*k:Τ���G�Wz��LѺ�",�b��&7�n�0��z��ër�.�w5u�n���`������@�@��qڅrg��U,�����˘~�4�o��y� ��H��UKZ������W7�{���;A��Jk�(��|;25it�����'��pj*/�����{���,��"�?� �&=w�b��R�Yox�:�|�K7'���M+�X��1YJ�x������k켬�����G,�k��O#R��[�0���}�HO�q��U+>���m(i��1�̻u���X��#�O���{i�([�8�p%a��J9��tT���U���
�#c��3�o?��L�BY6��Zε9W_=�����HZ8�*�nV�YR&�	n6�eO%d�gp�%������^5g���������N��D�x�>���l�]�	�q����Q���S��G9nz��d��8<ʛ���1Þ2.���q��0�Z�u($�0º��8�C�v���h�q�v)��%����Gsq�^(��d����[�}�z��1�QĄ�@��X_���
>��VLt�+@?㤒��?��X����K�ZyvQi���O�����CB������!>`��S��,�jA-W�B�6�-4� �$�l'��Z�C�O!��筳+�f�<�M1���ޕ����Ak�>T)�.|��Lo�R��X�b;�(ڱ>ꛋ�z�j:}�A$��rht>��j���7!�L���u�+�.��;Y���f��~GC!�����dܥ7Yܨ����N��-c53l@��uq�Q6��<�D
-N�m(���F�9퇊]D{>����X#@�%ԅ�����*v����yu)�#�K�$���~f۾N��qN0��Z��1�-��˓��q�J����.M���@M�VU&��Fp�v	s�+T�����TW9��>�slq�GP�DC<ۡ1E)<���HW�՞j�m�2}(?k|T*D#���	C�'�s�I~��Pvu.oz���3���.�*2o�����,-�خI���w���Չ|�F�^'K��r}�������j	o���8 
�2m<�$��F�.�U�z�&:C@�Af:_�L��˯I���y�����4SY��bV��~�(��%hR���Kz<�MSo�BvB���߇ڠ�"��R�5�J�_���W��e�^+�d���F�~ܙ<ϙpU�}�..����l*�P�.��Ji������jC+�Ō�9�᣺��5Mf��l���1?��+X��������k��c�/�f��)5��%L����΂�wPL�@�$Z� ����Ky��؉��8g�gD�'���me\�ak��A. ��X��)�8R� [�ѷ�+�W�P���oH ��b_1
���W�pR.��S�@�4o;�jS�^+w �R�{.�bnAZr�iRzo�rӦg�z^�)l�F�u�ʆN��9��_����]RKWT�A�y�cC�t.��#^��ڕ'&o����j4�s�T�CMG���0\k�,/�D&C� ��d��8S�b�"�H���_o�	�)f��@zB�t3`ƶ���6�O0����w/o�����s���/ʇjѳ�f�]K=h�μ�l�*���h@g��.17�W���ԵFHWc
��2P3Ѝ�����%�7ζ
��J���Mg��א�tu�>�\�������Q2�<*��b�����]�2�87��ѣ ��Ũ��f����ͤ�Ȕ�M��@5oX�C��K���fD� ���AO�Aޯ�+6���(�_�OZK��:�(���qQ%���g:Է�4��A����{�ό?\�ijj��$��ȧCieV�ScX����8�Ϟ��(����u��@��=���[�����{-_�TN�yW�4�k���F�Z��5T����6�	����XG!����b�H�.g�j�c�o�����+s~�H͆���"a���F��!��n�?4�U�%���gp�O�G�m���I������H�J����8+�$a/|�Ђ�%�#�U���%g���g!��^�6�'MuP��V9|��T�u�R-{�������������V�T��TӎLZZt�r#L��G� nG�5u)�" �I'���n�MC�1*��
V���ɋ��dw�nԓH��n�#���l\�����H=��&�3Nѭ�-�L����$s=;5���^."���U�A�aD�(ƕ���@\�5|�R�PãM��ט���*�}T�������P�-{��^Тe-Wty�,�
�W�Z9��i���>R�{\s(~�̀����B��гk�-�-%P��Qs�2�el �d.+k����r &����oSI��1D�h[�����`�5Il��/@�=�-�Yyc�K���=���݅�J	~1�w߬X@��w�e9�ā���z���@�TN
���~��ޯH�[��J�&�ƴ���!�a�7_�nÐ���sV�c����yx�f�Q"��^�l��e�1�/���u����ۋ,Z������z����k�\��TG��m�&�a���7����c�e=/NC-���־���S����R�(� �a�����m;i	2a���D+�Cp���ɀ�9��ĩ��m�(}�T= �cc��/	O�-t�`�1��NF�V9)�ߡ�>�g�9�m3چ6Hc_��שK�jYA�I\�2+ Ȍ6�2��6�V7����h��_���*W������*:��
.'/ht{�#��]���^�re�88��>���o5���ʨ�ɖʾ�X�����bZ�5a߇�����Y�� oi+�p�R"��E�Y�`+�ߞ��R����+H>���ې��W<g�I���\~������,Fp��*
B��5��y���1��lq�۶�<�;� ]H]�O���g	O8�GE�ą/���lq4/O���C�)��"��d.������b����������ss?��z�I�:��8��JdDtY�&P��������.�r蔪��]�}�/�l�c�n&�(�!�I[��b%�43��c�����������^���>����t��3���O��<8T�O��
aC��}W�M���'$�� ������x�5�<��˸��f���VџJ�V �t��?LFe�h��6kA p����@$T�%�I����D!�X	�T�Կ�e!���'Kuc��v\�3gx{V���P��!�9죀�,t��T�nJ�w9{<"���$5�{v��M��V?F��v��M��y�`t��m�������WC�|R�~w5���Ϝ���1�ɭի
[�3���[���t�2����H�6#���!s��תmF�v��x��s�oI�4`��[�p���p�w��?EXΦ_Ȫ�-U ��@J40E���ڢ����
|S�A��f~������#���p�>�ϙ�l�����i�����{4�e�Wl/� �k�#c���y�T����x��N��u�٪�<�ƀ|+{=S ��[���cKp���M�c"bp6(8��W&<������׼�W��F�m⍒�a��gc+�ՈiWc᭢Q��@�����F��\�u]<����03�/e������/�笿�uB�WS��3��އn�˴Ӳ�ߥ�~!�Y|����~͝y6'��(q�Dӝ$h
K�F��,q�?3=�AaNXCPc�l�Y�h��c^�~�f���8"*繗!rW�Nj���Nʸ�rwE'A��~�{��B����TP�� ψťZ���R2��z;@�,�7jc
���*Mî�z�}����y��I��o>�����/f���Ɛ�D>�G4�4C�XW~���ˠ���:a#��0$d&KyY�����sҝ��&��5L2�h7<!۔Fz��`�r���M4�pnt�>�F�]����2Î=V]�p��SDEDI�Vp��̌���Y"�o��'�N|oFZ��e�Y�G_-J�G���g�s.��TT���f>��2�`*��H��],�e?Gj_��f�.���0��K�E��☧��I�c]�L$�h�$�������9�j�G>YXrY�.��p�*R8�l.��g�밞��!u�ՉWj<�\�r� ��O�uhI�iż�@]{�=;ԘL��G'U~�V�?��rҿԍ|�wѬ�K�1�����5qFt���[2������uxQ���LEf3�GN#�#LN�T�ؒC��m�������Ǆ�>�B	iᇎ�PK8FAFc5{����ݠ��:��baX)o�_N����j��.Sŋj}��bȏ��eO�+(ӈ1�=�6wa�$%�ݍɖ�1��!xj}��|��5"�l���T,���<��_������F�����ک�oUU��'w��!���	�����B\gp�(�K�=�h�s���*�TE��9�Kb|�"�:֞��f.�n�_VN����\O�n��gG�'���㣀F%��)8��t���;b�+��|�J���{i���c�!6��?e_��]Ix7���$E=|�fw���+E���uu� *O����nS"vw8xp���?���e�NrG'�B�"�r���P��a��h�>-n�gsƩ�����yB��<�,Ҡ�F���T4p���U�	MM�ä�
�E;�6h�
�\p�KB�Z8��v+Gk�
�zK�ym��a���K�������Ͳ�JU��4)��ϑx&��¼��3d'M�y�τ�Q���?2�=��L@\9�U{
 �����~Ni=-D�6�e� ��8\L�YΊ�������J�d�lr:�oO-�+����Z6v���Q�����RV�6~�А�q�~g&��	����{�r�'�]g�:Ŷ�SC��3r%`�E��ѥq��'��U�R�̵�� ������$A�/�|����w�!af�$Ư��g����x^ ���7]:�&����0�����㯮m?6e�QƼ}���մ�*$��2T�;�ͨ69�����K��a���c���>Q*i7���ϐ�I���1ʗ{{�f��ci�& +�EP0�VTD�R��	��-�=8��)��N��h�&ھ�����2q�t�ds��V�,<��;*�e\�*���PG���e�P�O֯<���|�L���&pl���=R����@)S��D�a��(u�FX5���x��.%��f�ȪVS3�Wp� �U�M���r�n`�eu���'�ɖ`�d@�z���*�����7ñD�0:�6�O ݋A;����C�'z�땳і���/���u�m��+�N��U�5:A��0g����oV0�qyJ6{vn��Y�����+w焩��\#s�LW:L�,]���t^A�%3"ޫ��n⊷�8J��}6G,�mCa�,-��N4�j�l��1[l����[Yý4�(No;��z���&��EZ���;�E�t3�������_�Ct�=*1=M���~�J������>7�7D�xfJ���#��[g�80A,���'�w��W����y�)rl���=����F���n���}��m{���^AQ�X���~�	��U���>k��{{�`��Hr�M7EWJ���I��EsR
H{ �S��Lz��+���GdrN��f��QZ[��)�f;���H�$EK����5������~�a��kN	9��*�� ������b̓9x ���|ddr����Z*0m^�{WP1�aJ\R`�C���"rmѪ+$�p�F���}*L�#������=���� �8�q�����ݿ����.�=��w�R������=���ʮ�1�t�j��>����$J��w��(��fWV�[�	�q�j��z����4��x� "��P-7Y)��>���t\T�a�&]P��Lˀ����"	��т	�Z�
�\	��=HuvT��*'?��u}�"j8��%��
*Mb��)��Sz�?1;C�tP �{s˷���" ����\�Н�֔%���@�
'�S�����&�4�'i)���@��_$�1Cb�&j��C2�D4�yW���P�,��b�9�	��Ñ0��IͲ@�9$"���̉a����DЁl�����[ekb�ہs�U!�5&3Y�%�!5�B��t%�z�[��ۯ��é�J��Րz�Q�-�g��i���H}�>�v�wδI�Z�
����a�v�B@l����$�^�����[8�2��Ԫ't�������Q�`9��-��z�p�u��q�/c��e�q�~r��u�^���Z4��ޘ�8�EȧFLn�8��������{ۙ4h�p��%I`���<����C!�č�	���!]x��O�l�S�#L:�"�}�(섁h��f�B)�9^�j]�Ӑ8K#��N�@s�}��	�����ʙ2׆�O5��F��++I��Z3 ��hU�ah@eE�=}?y s`����x��Yi�)�K)�����,��gn�,�V8r���x�����se�^NҤ��.b��̀fy�w�Mg��^�7~�=�@�e�r/X��U����cSI/��ѿL ����q@�8�^C.Z��t�&y#QX�+��,+���X9j�Q*c���N�[#� �@yo�&")�D�_^A{�f>�+��@�90�zgV�h{V�n���	WXN�M�S�R��Eu>A�M0E�ӈhw���`�(�scƥ��ȃǤ۩B�D{-'H*�����K�w�&����,���[ʤ򁎩��.e�����t+-ǝ�m~��9>�Bm@�J9���S�I����)/CeWKC3�W\#�V��.s�VE�4Ѥt����zO��3����7�8����3I_�J�%@�	mX�c�������W��X}d��6����>�Rc�?���K�dU����F������8D� ��j�YL���5=�6�u�T�8v�R(���q$�/���_x����v��$��Dу�F�ڒ�z5b���L�!Mƹ��]�|p�
)�Y����Ȧ���-�6�1Xp�H�N�|�0�x_㭔�ƀ��2����C��O@���,R�W\�G��)Jx%�{,�̳n���ю5�����j�0���g�4��:�ʃ���'q�p=?`��)�6>gz���Y��b�v��Ŵ��&�����qI�,���_�7��s� �5�lI\U�ۈ#�[�iH-���5������u#��Ϗ~i�r�h�.�;�p�nЋ���S�ʲ�5
���)3Ύ�Nݝ����r��`�	V�:_i�f��z�2���Q!��hG��r����y 2V�j�&��۳�����&��	X�l��H�{|���Tay��u؀�!���*��b9j���S����@�ts�tI,��r_�yɆ#�6]�;�`����z�#��/P��╤�)߿�������K����X$w�l�O2M�!�W�R��fh���ҡ�[tQ�F�VD���nR�`.�qF��UL�?/�Ǯ#&HK�A��{�� ���R�N�	4ICI��\�K*�ε�3��a+%���o�O�h�#��Q Bڒ��6�-j��܎_��R��I�Ђ�Xp��6ܑ����5�N4�� i��~ևV��*��ݳO?���:������ �r���Uoo+	��y�dyGr��
����xF	i%l���L��C�,��\o(ְ�{�O��;kߐ�9�{A�%�4�@���"�!�s����L��>��7��q�E�F��}�5\�a}���S���#e(�W)���sA&��U'Ҳr����tߎ��%���2c��@<�X&/o6��<�~������T�<5]��0- Gd8|� ��*�Ѿ"�]C��-g7�n����v&����cMiDT^��x���P����{�1P��0��4�����[A���R(G��(�|f$��[���T���bd�sl؛0�*�#Dv9d�LXd�󁼍p�r���~'��??����Eo��_$�a.��`��G��j�l��PJI�p���Tprv	�v�mb��T��D3f�ǎ�U���"�z�>�5f���_>p��S�/�����&@ˁ<��l3Nțr���.���_	R��D~a|�&)��' ���|T��sJ�� �������b4��i�}��R�go|������N ���xW�qfy���\mvcD� e�}��0��7�o6��"H ��ġa�we�S��Պ��Pl��]�)���$�#��s�K@*Ze���{�Iv3�r¡2�D>ʍr������%4��A[c�Q���7�H� 7�b[�wu�ΐ0��k��k�޿+�)����֩:Vq��Ip�
�1,%}��nr#z2@#q�(^�pNڼ����_&��2��2~ɕ�v��>J-t3�j�9��$ۑ��} �9�F�M���=�Μ ���}ID4��#(8V�]�%���7�Kֶ�:����ZC�ֹUZ�'��eC�L<1�^ߋ��[�Fc�2����d~d�1)����P:��wEoH�mЈ��ce��^s3u���I��X�Q'(��`��n
�h�$��^� ���4���
[��c{^sD���_967aEك�B���P�[���[m�Hwƞ}��["�Y@b�Gl���z�a�(%'��Z	�W�(k�/y�("l�A�d�;v�7��n�;,�]������Ly{����TnZ�*-k��_3g�����t��b��X�uީ���pB+���h�xvSn[�r�B�O2�Ri)K�5-8{x��=��H@\V�ԡ㖻T{����\��*IV`߿v�$�g�ܧR�#��0��{R�J�Ra������zE�p�)H_�Wܸ*8�X��E5�����`�F�����C�����!2����;y�_�q{�������R�DS��0BcN]���^�x�~����MW�h�o���
pm&^��Tza|-�4c_$ewx�2�E��m�`��3f���\�fFTv��q���	B�j��$�u�q�ي��4�>dl_�1Gb���!;�\J**;PT_2@K��`݋��UR$��}�"^�!���`w�S�����V:����
'e��
9&jqy�*g�Ա��o�s�xV���5��J).�Z����(�)$��p���hA͵G�"��������y|[d�ݹЧϲ���7�[Vw(����ua\�7����1 9 Q~���X���MU��Դܽ���f��c����(�����Z������6bN��)�EO�����_�d{��C>/�a�JѨ�y�&�(�|�H""Y���#T�;������?uL.UzM�j�o|�؂�@�f�
`H[+}��]9�Q.�pl6�����$�C]g	Co��2�jk8|ޕr�j�L7�F@��yiQ�ےb�^??�ұ E�17�>�)o��F�nnn�m���;|4P����{ҽJ�rknmQ�x�������a_2	�Hj�i�;?FPAr�F�,~W�;���_��8VnBJ��]�i,�E�Ty���6��K�gLRGÆov�� �oJ�y=B��%�n�Fھ���Yx�o ���Y�'c���_�rf�� $!Tz���r�#G�b\/���	V�B��gx!����ڨ1<^"�(��֓��\E̼���Zj����1�������������w����;���}a�Ʌ"��s�4_(�Ъz(!̈t���K�M/\MF�j���<���:g�2{S�ǅ� /��	�΍���/k���	+/1��,./�?h�%�.��B1b��pR�x�����+w~��V�J��e��w/��5g͚�"8wv�A��xm/h�(Mi2ɕ��/ �;�=��\�rg�ٕ�g�M�Zd�Pޙ�4�f�;��D��@�j9X�T�/g 7��\�̏0>&�3=D��O�C��bop�Gf^'�h��0>J�t�a��wIp�T�S#����Ǟ|�C���%�nhXN��#�"h��R�}r}��?��s�8��~	�!�|b����1$�t���Np@���مk�0N ����]j�̅+m�I�(+^�b��V+Rs/�x�Y�Z����zN�zr�Fo|t���V���׳*�Ԩp�pѬ�mj=&�s��	TaLi��EČ�X��,�nVs�|�h�3������4��,g�l�I+����Y͉��>$?��o9zpWe;ok�m55Ǌ�� ���a�s��\������Q�Pn)A�148'�d�9��y�����䙨�ޓ���Ё-�AiL��r�s[̨�<:fGK%e���5�E=)�� ���6��^m�濃�`r�39#p�ꤋ����N+z��5@�����,8�PHRR�uG˳M'#�;�-�2���{�=���%f[��k{������0��[�.aavG2ܙRcM~v4���E�X��_o�7K���l$"��jy&��I\�Wz���pq�-
r�zw�ٶAy5���=�ޖv^d[��� �օ�1 �<�RCR�"[�_���@{hH�fy$d��-s-=�&t�ܴI��F%� v�ȥ6��r�$Io���Cě��J���y��-�Ü��m�+��,��Þ����y���EЮ��욒6s��9Nx�\o�_~ǆ(���<n�H��=�TL��ǁ�a�
UR?�}�i��Y��Ol�j��������+R�4TF'Z�t;Gm(��z�����7SmC�dP��b�/lh����eBi�Ԛ��G���>ο�l��<`�K�x�U�1�W����j9F_�<��=�E�A%Y�*�z
6-��H
�V�6'���+F��sVg�.��+K9��� }����O���Hp�X�W�Z�bK�\����q؍Y�י��%�f6he�
by��0R�]W�5MBP&������X�:/�j�͍�N�tי��<��R�TYB\�@�;S�j��Ϸ�YyBڑ4}B��[�q`�_�m?x>�\N�	'y�&����wJ	/`��}W������e��S�}�B�]����#�#D�������K�qrz �#���[���vZ�7�*��M?��9k�fd��n,f��?*��8ۋ�q��W l/����gފ���[%���fW��֝$(j�(��V3kT�+o0^�C�>�D���A����k��~ [Ed�������ב0f����;8���,2�͖��;�O����tE���3sC,��F�]:}���ߜd�L��[�Cf�6�F���Ls3?�� ������(�ΚU.溲�	�!�	�'�\��?G����g�����g<7VSB��`���}�W{/�x�SR�9�p������>.H?�oAH'���������93qYiǱ���	f�u2��̖O>* ͝Jµi�s��\�b:7�<�pg��3��"+�rvAfW�)7	�C �sj�dYc�V����I��ѐ]^"�J��(��PL`s*+|�#�F ��j�<<@RM��.W$�A���¶/��%��ӂ;�Ċ̊M!����hP��"('��ʷ��R��y��Z���2�h$pZ>�J
��:v���(���&������.WJi��$#DA2Mg��>�"�����X���\�N�j�H����`��{�m�B����b��
�0Πp�u;��`C3�9�))lo"���.�}Y�,��!����*s�s�1=���"�����yn@)ή���
���D�N�:a�9
c}q��)yl��k�'�L��Q ��G���bP#��"��y)��*ՠ��"��D�q�l���eb���dߖ���~
���,�8�B��]���D��Yi�Q7R��ܱ_���z�c��}��C���anC�����k�B/A�㔌��Ӕ��;�T����5#��؅|O.ͳ�qY����?z��F�Qo�v:���s[���F�P��[ �e����'�@G�f(J��+F״�'�S����+}`���n�Շ���vPY�9 =�l8�w6�w���������,����DVՐ� U����HΚc^�j�N�qc8Y�����4.�"+Yb��=i$��֢S�6�s���*2�^kkVؒ!*�h\��%��U�����e %�ʖ�@V )�_C�*�i����;���65�Ա���BO��_^r�ê���AJT(<)%��RS?�(G'"h�r�(��E!�A��&b�;0!�����{@����h����ʏ��t
T����?$��cP��#�D�7�4��Q�K``�j��+������Ƞ^�.���%��G�׀��},N-�&�?{�g!�83�tp ��dʜ9��J
��9�}�g *>�zv�s]�}H��2��2�Ѣ}T֮�am�yhL���x�YɁs�CHFi+��p�R�{A��/���^HsO��.��NGB�Pie��BO��\�J�s;�m j9�`�Y�%���Qq�۰[D�[uK�b��	���<� ���#%�;��UXΆT��W���b�ӂ^/�;�4���Z)�c�QN߅]2+�
i*%�a��q����']T�ba����!s��#^b鬾ZHR�nD����k�(��<��F2iԊ���s�����ux�6�\�1�����G�*0w���nhb����}p>�IPa$FN��f=��ZSf^�S�s���i�����SfFʃ���'I<�[Z����]���2׬��zW�[�CԷ�+AUګ׆��@�e
tܳ��-ߘMn9�MN���%�'�u�<�,�_%�rQ:0q�A�.s�3�����a+�=��V�z�g�x��kh�.��H;�|���u:��H��j��I�����v�Ufj;	}-��IU#K{S��ƟK%������򒎹�1Q��=q��T��"ga� �K�� WM���	�.S����Gar>�*�fW��%�o����Ϻ�;�*�0��D��x��	ڀ8�/p�	UX	�(O���[b��������ѣ���Ͽ��I= ��~j�����[��]���.0&��"�$��[z�x�G;�$�*���ƼSU�jING-%����R�:w	�])a�.&>�e0���T"\?��g�V��B'�G)�$>�x[HXq4�x��;��>ܟ�'��"����:�c����x#�<���Z]����Y��>'����IJ��0W�'����1d-�.����1��"nrތ�g�ʊX>��Sdj��=
����z|3�X��M���g�g=|�Z��=ɗJ�sՇ0��5?�� ^�?@Y��?�KB5m�2"_�+��$����չ3�� =�h��_|ֵ��Q�>z��jo5̔�I�Xh�p�����?�<��R�S�S�y��}/�I�4HT�y+���Ԡ,��'��3�=ƀd��^�0�̎�����֘mml��tj��պ���r~B6�B�˨zϟ�	/�EKP���5���@�i%�$|�#y�۽�������(M�O':srq����pN�ɪ6�(/�x-��5��5�&t��RT�gJ�y�VIt��edij��ML|�[k����;�#]U4h�-]N�(�Gĭ��'�����K|��35|�`��<ᣩ��7v�Y*��,IKAX_=8�tǹƛ5��1���y�[�	����i�)5�tM�eMP�i�bB]��O��S	O�7�s�v��N��	!z��^�إO����Bט0�=���h����5�]T�hK_B:�t˛!���a���_������v��x�Q�
A3o[D�:�`����j�+"�{PCNlr���[��rp�	 ��7v�3�|�7���Aw�A�,�!۳}l;0rׄ������Z�+�hs[��+����)��d<!�2�a��>��Y�d�A���xb =X���nO��F�gJ@��,
��|H2Sq�(Eز7����}�D�?���J8wo��IC?��*���'v��-�F|�˦�Z���Ӝ���y7�ʄR�<��|�L6���u�6���ѥ�Q�/���Yi|���y���8$
|�{��7��h�ґ�j"�����J�鞄
r,� ���0�󣛓$��M�U�K����*w��e %�۹���>}�E-Ҕ"kD��!5&iЎ}�Mi�$שc��7+��^<�D�I6dߑGa/� ��gs��?�_}�9z&�8�5�,�i�t��=�&L�A��hܠͣ���FR,����;G��r��|���؏FP���ۤV�ʫ�l�v"��C�ʪ��K1����!"&C>..�Td,�5�<�XS�z3�V��26�*� G��h��J\����s�;��t�� =�"-
V5q��㺳*�e�|���2�]�k�B�x���܀�A�Yg5�x�M4!1�@F����V J{t��Q�s#BQs'��st)Nw����^��\��c��|e�Bwј0�,���h�3����Xڷ���	�������?�vep�~�ʙ3D�ND�Z�� �������Y�v�]��\qx.?�)����4*�����D��y�F����]�f�� (^IT%MGHğT���ўod�UI�P��/���)Va���n%�a�%�CPR&��h�2|�ͷ��*O�����@:� ]�s���x���������vʠ(�)�����l`�fa3�Y��kT��@���A���OL����A"r�^am9}����i|����ʡ%y���d�H^Tm���o�π7��N���s�h�����+:�����t�[�W����G/��J*'��	�X w�����bCFbw�8NEZ��* p�t���	0�����	32��N^��h��bH��'Cl�|E��8��@��R<��� *�~E�tY�l<�U@��THQ�z^¹J�^E6*$r!ݛ��`cg9�7�K�1���gof�+��x^��T�K���4ał�r���̍N!!\�q�s��K�f��^��:b�*��<���kG�1���CUb���S����f
�y��Ew��u�U�4���E�pO I�4�ʰ�R,1�`�ѾVj��&�4i���;��vԊ�8;�Gk�:m��=���H�#���44��Ί�=-JF�Ox���һ�%w�{v����·3u���քQ�k���5��{d
I��#��gB��x��LŎ��.O.��$d�"�g�&����FE];F˹��#m,B��37uc`���mWL������ �������f�G`�f�'��E| ����g*$��e��$gc��i�j4�E�������t�U�N��A����HE�Ι^6)�б�=C�Ĥ�I��d�#��fn�)���ꪥD4�"/%Rm>�;߽b���פN����BD��ȼ�}�:��?9|��x��?1�;ݎ�Z��J�O ��G��]kY��bu�y��A���*��x�/o���T�[��V��kp=".���N� �d���lLa�Xp�����:����d�� �tL�<7��⇽T/�Y���
r�.�K呉�
�r���M����� �r����B���EO��n0v,�)ޤS�|]�-��OV�M��z5�Q�e;���/%�Y�ze&��4�z��g���{#
�_���� �VZ~�Z�Mk,�Yz4���.����:��k�S�`�a�c<�����r5��6�$j7)"u�|94�w�l2�$5���83�h@|�tҒ�'۹�8Kg�� _^L��g/4O!v_�����pel�(TA�fGٴ]m/3���e�%���4]|�؍��˾��Pg�ɯ-����,�ǰL$��/�&d-�G��أ|cǄ�e�qҦ�Ћ�|��E:�,����mÛ|0caׁ��rO!��Y�H(S��ZD6����ސ��s���&��~�MO�:�L��.քw��A�kM�mԑ�m
�����CKӆ�AC��?~�ഗE���YQ��|5�׋��;d�u�[��o����d��7��y�=''4H���$�H���:��o{���VTț��T��>�EGu�>�c�v+9���<m�O�m��[�:oQƯo���Kw�"[����v*���������l�h����5�%X�e����S�嶽㇯�[N�W0�*P9�k��	30�(���l�s�(�4��Vcqj�	\��f@0���$~�v��M7Ϊ4�>�'fd#t2�"�=��n�1Ȃ�fƮUM���!���!b��a���f�����"c1͙:K���9��[�S����"MqE��̑�&�g�]YT���{��~��O&o_��M�M��C�Α��������c,i��!>[N��9뙄����Jd%�{0�AhK�jED1$��i�p;��{$�I�U�}:[�M�Y����c|�uhf��O�#��ɝӠ�\���2��BX�%8t-F�T&m0D��7�gz�T�9�˩H����ߝ]���3��t?�Íҵ��$5�P����m�(���R�[0{2{Cޯ�ꭶ�ʄ=n4ݮ8w9~چ��!���[�*��1���Ew.!�vc�^���ۂ-n�5i]�T9�C��Ū�l�����I(�̏G�p��6�V��2�r�g
>;�i����d�y>�^t�a�QG �
�U�Cl:Z/�� H������i!�/��!�[���/u�E���
�w�����9�����LZ :�Q���;B��U�m�d���HI�ъ���w���^�K��	̛�\l�$<����#z���~w*f��8�L��6$�.��7j��m��s]���)CjV--����t�v65�/�Kz��mY��+�\�C��� 	��ml�����V���x���Ny׶�j*}�vn.����{=��q��d�ԗ �p"/^�6�w�My�qK�>�b
� ^0�ɿ����0yhy��M��s�-�&N1fN���]/��c���i�=��e�$S~��Uc2�,7>%�NL�-��M^�;@�V�&��f�J("�m��^FW�_��)r7R��Ņ��3���</3 �J������Ԭek�r�앣���|�b'�<'a]]��C=vGI�a���h��q-���B�� �+��,�uՀ@�#C��v%�Θ�r�BQ��3m�(���P�Ola�˲+��2$U��dK��mf�[�XS�h�+��7�ߞ�x��m�ME'��!�h��ʋҦU�d'<���jҬ�
Aԝ������j�l�`�����T{K�c�^4�`5��b��x���~.�P� ���yw����Y�h�F/��0��df�5�Z��
�R5N����W �W�_�4R�V�>_�����5w�����UP���Y�!��̲��Wtd` S�y�!��5��&*���C�l�����v���&ڪGc����dI��w檹q�b���J���k�͒���b�: �l>ڹ'��1Iw��{{�q�!(䕖K��'`'4�k�T<x�$Q'D_�����:��^� 0"O�GAhV�����2�t^�8W�_�r�պ��T���U�����d���R|��hK�X<n�A��K��q��W��x�eMM��t����˜ú��Ӧ�Η�}ωϓۇ���h�z	>g2"��v����m x��E}	�R
[��iN���*�Qtl�X2A�&=J�'���[f��k�E������������>0�k���lJv� D���j�It����J�(��s`�bo������	ڠ}�,r�����:7	E0�dK��<��<�)�m\��w�-3z�����IN�P��c�ל	���� ��S%�A�%\�"�;d�Ik��,Z�KlvI�ĸO|�ki���cv6�����3�b�&+�J�
�#/�LG�c����0�`�}M;��I*��g�#s�`��ijD&��4�F�{Np�x%Lf�6�|��#��p!/?a��H����n�A�f�1x�c\���Fɻ�d��ceQ(cqghQ-kӓ�@�U�.X;��su<c��	~v��J��7�E�@i�g�EO�+��˾q���H��Ym+�o�g�~�<� As3L�-v��bL0����[ܫ��Hޓ�t���T����|-��½�H �je0�rD����<B�R̸I�v��nK��}É���+o
8�3�]�h�ʲ�oqu��@)T��`�LFƆ��c���V�ʔ&�P�|?��e��\�Ī 妣����9��uO��C��W
j�n:!\V%��Sf~��d&(���c�V��&�#�p ��#�3R�}^�>^p��,�W�1�Ѱ�h��v�,�F��ۍ�U-����5�0�:?(�i�!�jm:�3U7*�CT(�[Z%�`���&	ښՂ��ӑ�<�����E���N�rz�b֠���owח��°�al�ìW;�G��������?�+��j�N �g��ڌXYy� Z�t �i�'|��������� 1����I��/В:�t�#��B�� �G��pGQv����H���m�w%u�}�@��kgm���z�+���t�u�ab_�N0�%O�Y����><<m���d{p(�#Y��2�������w��^^U剋�����,�A�6�=�խFmo5�I����~ɨ�|c�	��h�%q���,X����J�g��{�&E��b��=�}�I@!�?5��2��n� u�HO��1N�����x���&�-��aR�˛.��&@3`=!
���̅u��񢨇�r`��I��,��!D�d�;�s�e� �F��H�8<������~��*ӯ����5���G'S��:*9�����3�53� 8J�a���F�k68+"�n[��lu�x���?`����$���	�KƓ�֊��ݑE������'��g}0l� ����nj���v���;,�9BVi� y��m$���C�����Sߨ~����S^v	���+iT����Ǚ�!r�K;��N-G�XryLf�Q&�`���%��-ƴ��� �3�?���k|�9�&�9�A��Ɍ�()�y�1vI��-|
�=�ި�٢�$z=,����m?D#>��Z�����F\&� ��ӵ�խ����,l��B,���bXs�K��ţƞ��B�L�䗲�x1]_BP��>��_�մ�=2x8I�~5@�~�9]��e�)gq�%+!��JҞ��w[X��� .��tw?5O��8�q#^`��B{�ì~�vA�.6 -8hou��>��A��x��ܽ��Q���PO5B�9o��[f q}*vI5�R�
 Ƹj����R4�pә�h���J�:����;���_^�F������H���ލ2J���f�� D#>�(j�."I��b�ꇹ�]�o���q���l+����g�( ������P�Q�5�X�ќZN1S4�«SvP�ngsf��h�Ɖ�ڤr�2�K5p��v�y��C�G���u��9=Y5��+��֭�6/u]�2q���%^ߍ�ї+fj�H���Y��x�o&n�ȑm���͢�2��^MO����B(`��+���Fy"<��G#
��gOA��G��$�Oc~�ak�7;|�kKg-�,+��w`�{y�含@������f Bc�v��I@��e�-.�3__�����C�?nJ�1ph�ڿ�#@R9'M�3��rM��1;�B�쎮r���,�d~��7� ���J�F�Rѻ�gK*CFt'��3��7��z�@�?����~'���\�wd�-��g ��B�(���>n4���I�%`M�Łz��_�\�ʣa�
���!������.O$��e�Lt�vq+(����HD���00Z�gCw-_���UaE�k%�@SjT�
9ƌ�"u?s�WV܈�h�חo�}C2�(&v�b-H/�O6�-�S�U^�G�}��DH7�b��F���h}��u"x�SW�����;[@�DD��	p#�*�p-Nc���!����8%Ӹ�Z�,.*��e s
�3إ��%#û����郏��m�ye�������k
p�%��t�w�)�@��c.Z�GD�����7K���~���t��^�'R�����ｨHa��Te�St�����5��]@s*NQ�AlS"��LB�4�Mz6Ȍ�O��h
4��SqDV_`�a��,u��Od���u6)��x�l�W��#Z3'��"�����4Q�<���ư�=Kt������t�U�yc��5�+^)\1ߐ팆/�&ୡaz�W�_��q���I�����B���[�h,��$qz��
��v)�����l����vL���3�U�p��DB���	CW���3a�2~&���c�pq�����P��h<�i��c,ds��w����^�����:�BÓ8Ȋ�?x5�g�<ɷt�\5u��ߩ/.,�(Ȁ��Tl�+�e�HV��.,c #i�GB�fl�8�2W�
)Vq��l����z���5'1W��V�R�m!�ɏ�r���}�u����%�J��
/��J[���|��X�,�w]����=]F�V���� �:n���gye�r��6%����Y����f���= ��C<oSʗ5ږ!o:TUp��P�c~��a��J6%�<e��P�n�0v�չΒ��v��0�(�f<��FĶD�HoJ�T݋"��.2ݟ�>.��C�"ߊ�n��_~gE�<3�SW��O����L�k5��p��iqVXu<� ��:�x5�+�wÈ��X���-�_T������$��xp-O�G� �Ӝ�C���Еg7"�W��]��(�QC9C]cxAD�P@�R�cx�g�A�v��C	��}mI�!�F�渭�o��C~I��ٯF����ő!�˱����d��6=52���}����Ԉ���a�qm5�*�⨒e��̷�Scf�뭤�)�(=��V�����c�{CÞtF��&�E�!p��'1��Cu���8�G��m���T��� ����Z�I���#��d�A��3K�!�w��7Y�\��<�ҍY+y�9Ra��_��� ��`.��z"��#ܺ��rSC/�����~ua-�����#*�T������Cç)���&K���!�-��:�����z�q�bMyb��C�ُ�����/�LT�8V�J���@r���$0/}��L��e��l�{���)/o�@�#&�Ӓp���X���"g~�1��}x[K�xs6��`�굳뾷���Sp�Yof`O�AA;*�����2��8����&� ?�L{�������[��]�#$T�Z�<�o>qEC�8x�"�Ũ_rq����b�̆3�!��:�n�=�b^ sj&����!稫��}cJ� �s�T8��g�tr���^�=K���\K�-�5t'J������К���F0����난�+T����<�ZQ�
��t����R���]�������������ЫQWU��=��ި�T�0K�X��T��	#����fX��)}���pO�'tp�	��c���D:\E6�l�F���DGi���.�ž�!� ��2p�2�ӑLd���Z��bd���G��fHDc��=:�J����*b�ѥ�� *�W[���`�xU����n����'&Mb@9�vF�K��.�#G�BV����r�x�C]�GU�EgG�x
3��r�-�c}5ր���K1|�~�/!��4Dﶹ>a7QT̛��i���c(s^	1´W1�8���G3��,�,�k7@�C���� Vn��b#�d�+QX|�L���B4�h/��~�����|8�WL풳ĳ��'Q�8d�����W�Q�F �H�7�?/��6�{�$ٙ��oB��送�a��Zyu�N~_�ߒ�K :�W��(w���/���X���W9����p �D�ܧ2�6�DJ��%��z�L6�E��A��S�g�>�q�bA(��k,2g�fS��I�V+K��v���9�90U�˖ ;����*̗�.�H���ư�ǀ~f ���;�E�K$�:ª�͓��B}��.y�Őd5Vs�E�.�uG&;L��ODj�������v�K(��3k�>��N�uSO�is�U_�j�tp���m�c���06'���<e���]����(���X6	���z���H�q}�c?�4@��L�<��Q�+��4�c��sH?���1���Z�ôˏG�@�.�� 5��m��J�kk�*e�]G�.X7.a�mk�Z��g�֯/����^`�b�3mS_T�"���m�M��(&��$�����3G�w�=i���&g�Y����&��O���5W)���O����o^Q����e��BL��7?@�C���aI7�k�4��s�aW�x�[E!�3�ꊘ�nUϯ�� ;����f~T��؊t����4o�L���jarN�¨.����i1 ����E��!1��
}�إw����j*��J�s 
a<A�z�7５��4�P�S�s��;�]Z���]́��e&�"��&��=\[. 13Ox���C�b�t%M�,�:�V�}|ޜ���Y�qpx��F9�� k��N���`��tseO;;�cZM�-�E�?�����A!�\���y`�:O�t���r^%���xjG�|��ŀ*3DLR��m���v&��C�TYQ���0���0��Ԩ��4ӡ�}5?�y����j�uv}	a6݋V�����V���K��ƭ9��Z~څ�g��	��2�9U>��x��T^��1�O�t4�E��#"Q�����.X����[����	fK��n�!�jK=*�Jv��[����k�]d����t
/
I���!pR*�)�z^~)V}ᷲu"��dy�r���{���2��g�w ���ڍ��@��2#΅O}sV=�6�9�u5�+SLW�k��\M��v��<��򓉉���W���B��"8(���&��������x����G���}ۃ����<������d�^���C�|�_1~ 3�6��p��Ƙ봎�b���.���dv��
P���ץ"Y��-Mo< ��ݵD�y�H��_b+�K`�rs�␑��= �M��v��w�8��l��D�R>��|�\�o6L�S]�2R���S����A�c0	۝#5٪э�,e0OJ� ��Ҋ�KB�v���)�gR��f��R��@��K\�{,��Z���%CJ*v�	YӜw��F� 4��?�^�Citp���Rc�9G={��0�wi���_ME�]��$k�A%@��ps]։� ��oa᪵yd�����.a1�5�tݤu�����;~���an��/�û����=���LT���&.�xzÙlJR�Ɇ��� ���2�S��ƪ:nȓBaB3��E�����c�ȟ� �v�֑g���`Qf��� gز���zS,N ���H��'1�u�W G;���f̮e���tø@]��V�J�o��F�~�C�|7FU�U�(�}ڂpwN��UY��I�݊�����&���ծA)tom���6N?䪸CJ�Nt<������b��iN���%��J�0��9#f'nZ����Iô�h�:� 9��"�&�q����8�~�f���;��T�syt��1��:ɬf8�H�_ݘ7N`t�����s�5�_���������")�� ]��7ڍ�P��DY��;t�un�Xt>ܟŧ��*K:�?�`��!T�2���_�.l�2��E6��:�B��)%8!)n����B �*�9DC�-i�N�,��l�4J5'�ꋀ5�H����v�dϒ�T�{h��)d�~%7ֻ�9n}�\�Bڂ��r�F�����~F|i�j�	6-C5K���(t��ݕ/g�A���L�Fa	�{���/o(	S������	2���+�c1�J9m ��d�����)��4�3@�EE�\׷n�q�s`_�w��8�~�c,�1,�b(���\�#m�@ɘ�8wY�|QO�����4X�و`X~@v��Z&%�l�T� ˇ����Ush����~��5���OfIؓ� {"S�L�zX��@Lة^9���^��2:nT�cj��K��Y�����E�z,���k��0���f-��U��О�J�d���̸�`��bR���؊i }5˜󴥂���eH߆\���vP�+��-Cy��Hֵ0�\)��'Be�{��E���(������-�	�U��u��i�ѿ7T����D5A�ڶ� � GF��B���Y���.][z�bŗ?S���F1	��(I=������H�''�KE ����aM�f�i\���`�=��Ej\���1U}E5�,�1�|3j�?+�ZB��T�\�!�]�z�I��ߺ�z�H�SU��֘{g�sV�%�a�z���Z��W�B*6~:���6뿝�	��L"���_��q;�^5��.�%���wt5o��>t~#��z��̈.幊f]���'I��!�/���P=��u�����@`�?�IG�c~�j'�4�3��NF+�Y��!�+&�%�[X��K�P#j�F�d}��J����r4�Mdx������I�t���(v-}�v����x��W^�bŋz~�U�>c����W4�s�q<*'�=�kO��������5�������vW){��Q'�d?QX-��p@���i�=&��@E��v�U�����ʼ��Ly�:ܔ��竏�x��������}?`;/�*��{⌀��� �?��pE����������>H���_��r��c��߹��_��:+�0d�q��S^kT��"�y����!�m�eE���3mp�ղ4������JbwI��0>��"v#.������6����C�hR3M.n)��ʅ]�]����t}aev����i�[�]3q�D�S  �zQ�d��Tʉ;bj	_{��3	55�dN���<Y����@S�'��`�'�fv5�+��U4!F�Ο̙�T$��Q���z1 E����t��]s�c��Vg+B���N�H����A�Z��1��+��M���u��E���+;���� a��
𗇝٬g�v���f���0���;%9KZ�F�V���+����<��9� ��;st��Ө�hPX��p���������E�D!�7���Mq��"���oE����Q���	T��f%d)v5&���ȯ��M����x���d�67�iM���	;yT������c5�o��<�b
���ޙ�3�,9ln�"�f�I��oz��,$��?9@��=�������W�� �U ���ٚI�����j�_�I���-����J���HW�U|��G@�6g(�fJB
&����?"�2�Uy�x.E�X��g��!$R���d��C���h���@%��q4���[Sc:2������sOh��S����}�L �=v���C�O���~�`Í����L�xG����mP�_�<�;-��Z�;DWl
�Ήt��FAU�9�ſ�{
�or��ONh0�/A�Pb1y6U-�vH��p��*�T�v[���ģ��Q�q�9��H�|��!�*ۜ�I�h��[#G���f��.���s�3=H8�|�/�}zXLh7U$D/
�ԥ �M�S�=B���V�8�D[��d��ѫ�`�e�&P�Y���f�{�wZ�7�)cɂ������6:&��6��>o{�mI)p�̹���|���0��f�jj]rf�s�7�A��YK��#��);W�y�0��)��V�(��c����L�A�.��Ǌl��J;�y�1�N- OER�S��T�_�b`��6,,��~�P�V���5N��
�݅t�u�NX�#9�:�I�ݥ:�_��C���X�+�mWu�	%���=N����z�c6�N�I���7)'E�A�l�+ٸ4~-�@����.cn\�ȏmB���͇�>֩�d"�s:���Su�K�g�#���<��dv�5ѩf.���C.�h#���Գ��߃��.aǄ���J%�{L����Xc.��C�٥��.�C^v��QSjk@��^�Y�F@��M��WA���J��� ��Q"�G5&-$͢;��0_��u�Xy���[�q�Kd8�)@k���bh��.Fq/�
I5l���`�v -H@B�D��3��i�g9l�"�Q�`m~ ~���7uʩc.B�[7��<���("k0��hܲ��Ii��_ �E��*o�r���0�/���X�kͅ_��C+rQ�B2<��0���Ҭ�M(\�J����u��_?�"�j�F�h*���[s� iI!E���%Um@*�n��ҷ���oz�V22�#'�^qb% �[}gz� �s�L,�\���:���8+�ڍ����A,����;3���G����k��Y)�Q�'Fh~��H��ۯ���G��������Rb�[�Eg�c%� M���y0��s�9ZO����·&�����{���4�/�\��U�+�� �e��5��D��t͇ۡ�����5d��ڒ����l儱�<M����ʞ�D���γ�/������J4��9޴�9��3�����X�5�9y�LM/r�[E<�@��LI��)+���P1���K�8pe�`Dat���u�`��v�C�A���Pʱ�(h0����y��5%���>g����N���I�l LT"�VH��P@�a7���ט�2T����@*1?9�V�۞X�.������*eM��k���6C_�0��W��o�r�-����H���<t���B|����}��r�����R�7H҈k��3Z�F`���M���%E$�6Ȧ���֞�N*�N`F�MR�낍����t.�wtc��E�?�2��:�I�����	��&#��:��Ɠ]���ң˙����*C�+�8w��}��f��QU��8[?|G6U.̴;�m�f
錝�y�ɓ�z�㔹�pF�v)?N���ONb��_0�f���[��wT�m2�e S��������A���F���Ks�˔`�EM	FW�~?�g�Wy�-�gYdC&mS�)W�'�����gI*]�Gab�a��O�򪢂�f~���}����K�8!p������b�I�ej��;8�Z�������Q�MJ��?.��p���GJiB��J�y~%@�g3�����k1�Q�m��ҵ��9㴊C�����JO�?�(5wW~�zB�4jz0 kE�闲&l��v��3H���'�RH��qǽ8O����o`)��x��>>~��](5-�Q΁�5r�V��O��ޱ�x� }�2�<��_j��b�S`:S�^U���)p�Lot�s�.�	X���B��4�A����{��Γ��d�֚���;���J��E��y`��9@��%��Иű@O�Rƹ�
�%t�R 
-vV�q�B,�.fDT}V�Jy[J�1�A��S�$k�蓾��t�ծ<toh��'��Vj��C{Q���1��;�{��i/��GM>DgcH D{�,��fA<��� Fʉ*���.�r�t�za �"�%l*R�ζ�X�_]�M��#����9�f�	h��{�,�p�Õ�J���_s�s��l���i�ƦVw\2�����z�-�ݚu{kN�F�Z�8��(b���C#��"��M�r7��o�Y.�MHG^vo9��
�:bT;�x:W��d �L�&�FT����a�^N�F@�e&օP�Vt������ɐ�	��g��[6�٥X����q��XK��'��Z6v��K�~!�P�b��{�+&��s�]>�Z0u;b�ZO��jѼ�DZ��	v�߰��U���5O`�V/-��56���L�0N������\�e�.��AￌP?F_Vٞ��3��Z����@���2�����l���F��ǯFp�3}�A�khsgY�<d�3	��z���c����ꇷ��hq���\y�GIy1��f�JZ�4����(+���Y�e}�14�&ei͛����gIcЁo#8M�{۽Ɛ��H$����S�$��������@M�?�	�a̝���:|}�E%��Jk���2�MH\L��s���__�y}V̈�ݓ�=HQ�f�F~\�>g�����/Y�Mo�QiY�����?���zj��V�y��+�pg+u&ߌ x��t������.N�[ʴ!Ee��Z�p<����}d����|a8�����3�Uⷩ���]fT��wu]�O�0��]i�v��T(�5���1�8�&�bd��.>�Hw�{\Sd�W���m�SM�|g�T�~�͞���!R�������q��Pz,n�$�{�<ȕ��"@� b�\2�o�B��du6x�Y�W��s27a�m��*�HmVH��K°߱�e;o�CH�˚?|b�s��cd(���hO���*��M����U���.�'R`�~5MЖ������W�~�:�
��=��l
�@�|�0Ǩ$�a��y)����_���m�*9b�R\�Z�*7��/�s������Ps�m\V� �e6�5����2�_�$y�V4sT?���pх�Pg�Z��M5 c��W�R�Ε=�Y� ӒD}���n���3h�S++r�����"|�����q���ӎb@��������<�*'�����ut���� 9�!�Og��m[yp�� ����떕L���I�A��Ss�w>��_���T�P�o��[鉰�݆��
� EjǤ��_k#T��[e�2
h�r�P�[�D�{�1vӮ�/G�-��Z,z��L1�29>�-r	�q����2�W�/d<���z!�X���3��ל<�1��W���U;��Y�	;r�Yk����%|a�����c�p���x��Wm��[�v�b�92d�;* ��s6z�vsbi,��	c6.�B�}��۾	���寮�cH{5x�^oA-�4�*�Wo��px_ߟ�@�]S4��%9�S�@l�)�[��~>�����
㽃^�sН_�>��2k�`Q�9Y��6�ٝG9q̘BǼrP�[B�f^?&�B90�u:J�6-���<�rSL���l:93"s�ZR��4�ܫ���0؀A��Й�3!�03b�q@_\��޵�A�\1carf��l�F�~m(60�S��#�?�P��	�%%t�.�9X��gD�=M.l4r���CXW#�ay�_)2�P����p.^v�`�~+�q>|�a���ظ1�r��G�_=�T��̩��r��r���3��N+��J�zhO,�_�bk3ŕ�U"Ajg��_�0UHm5����H`�;pq�\�J4m֫Ix"�"E���t(������cb�k����Ga��ؙ���-�~�n�s�L�'��P�z<����\���t˒���V�<_^_Z������p��՚��%/9y)�k�%Y�d�D��;�Z��������%ӦE�?C;C�>bTy;e#U�7��nl#B�(��9ȶEK�^+p��C���s��O|�����+5촿!/�rV��G�֙Dq�1�ו�P���ة��/Rz�teG�!<�t\#�<�j�:��M�-TuP� �q�%�ݗ��۩�e}�������n���᭡�K-M6�J�Zck�9I
�a���ػqg�zP�U?\�iM�&�]Y�����$��W7 �H~��i�$�M�}4��#I^A�UE&�A%	���׆�Sv�Ʉ4��K�3�ѥ-tBW>��E|�t�m8�,��ǿ�`�#z��w�ھ(7.1Z��Uguw%J`��c-�t��~�xJ[���~B����
7�rܖ��$����HU��̻F�&ڼ	��[v�ƂK�`Ş�B�ܞ��n�y]����Dy��v<<��鞘  f�ᚥ�h�5���#o�:^Ȱ�5�����]�V��`�Ff$��%��y��i�S���:���� _d��o���DC�сq��Y3G���k����x�rµ��8�bz���kD�yNP���rI����J�/�s�*��� N�p�^.&k�A�ȽS�.�t�$[s�H��N��晓7�~('+�Z9C���fw��9��~�_6}N�객q����cm$�5s���N%X���{������n&ɘ\�d!������_�?ah<�c��>���G��KO1�b^-H|�K�:��8f6۬�~���V�ֳ!Y�/��13l�nU����4/�M�2���Ÿ��x�ӯ������IK3�� M�M}+Cq�^0$s� �=���	^5Bȧ� ��y�)�� �&��-f���.�Mo�I�}���ec��L���\螛*Fy7��Gq��=�r\`T����-�s�k>_�^.ڷ"R>`�!�<D�8�%�+�����n���g�y�����h�L�<Y��봚.΋̬�2%G�������	��6��`7���R�Ϣ�[���|�o���K cX��t�^^���k���|P�.�z��]��04����/"��p���#�Z���<ɑH��tᣏ0��+�,q����N3�-^� y��)�b�L
b">&��Q�?+���Т���u	هw�!z�c�Zj�0/�jݿk��f�]�����1�ņ��>���rŰ��Ķ8�T`����YL��$R�o(�f8��*�V.�1���((9�9� ��J=FP��lZv�SCZ�ϵ&�n�����Џ�?��_+���W� ���(�+a���Go�o4L�c�`�a����J�w�0=��=��_�̷ ����}ɐ#�������{����6Kl����<%9����җk�\�|�Z�[�zC���M!,],�â�̊R#� �m��!w���b=��pk�7���.���Em��!qT;{�Ǿ���,HHl��@��K�^V�Y]��jIu*~�(���	t�^�	�+=������X�!b��8l��رw���{� ĺ�"�-�����7.�P�̻��j.���aЂ[�c[�2�E)n�^m��;�ț&�<���4�b���`(t�"`PO���Tl6˧"q���0�!$�e�nv��	�������jM�vD� �*��ő�����PXWo&4�kԡ�pdc(�t.�'�u�(.҄RK�4e�	�[�nl�0���_ߵV^�N�d ���I4�p�d�Em.�i���<�؄ڸ$#
L��o���8��p��|��I�����yst��/C��Xkubq��で��С".$u�郷'R@�'�����j.A�b�Ob��`�co��e���J*��󯈦]�2��"������O~l���AVr9��q�iCI"w{t��2#���m9]zjQRr����U�ZK��s+p^�:�AfY�k��?�T��6�6
��#q_:�(ۉ�u}{&�7��;ܟ�F����/�Ye������T:���qF��Z⻮�	�jɋ=	��B��7��7�5]��#&�)���QMB|��瑒rXE�������L2Gm�2��f��laP�ɧ-P���/Y5���������3�K�Gh�*Y?��`�P���w���č��%��}f��j���/���%���W�jK�j��f{O\U����,9���k��ٴ�}�`�_/4l����x)5���h�/#�>���(��m���*\���k����+u$�fQ~��ABA�k��'z@b)O�^C����
�P<w���F9 Z^j�Z^ԥ�PJ|�U}P����Cg	��a�G����^�4�̆�N���X��f'����Sju��� -|o�	ģX'k�m�:�o���'�D�1 �h���?��Q� ��X����p\:�}GH��)������"������V��Df=ODqC�b������c���ku|�ɱ
���K��G4�����;	z�`S�>g���{j��	g���K��zHYT��� �Sc#�Cj��2�����;��_h��.F�6��2;t�B��g��:;u��j5�*Ts�av���Rr�����Rj�������"�o/I�?�R;�h����D�&dfL�Qz�\r�2�`Ln���qRQ$wvS�p��_@����
'*yt @x���u@�3Z��<@��nX�"�绸"|����T��ո����e�94��⬣y�Pn�pr��N?\�8�_Ɯ�]Ww
�=��#Tx�N�Xhh6�|�o�w-:9_��������_��r1�3�t�9��~�Q��߭ hr�{[j�ޞi'�6!�1?*%1�k�Y"�ӥ H�h)f�6����vv\ص7�g��U��U�p��5HA�Ϸ28By+C�E��B��B�^?�Zyh��"ӗ�&�VpV�����L���׺�Z����p�!Yl!{2c�	�LM_��}�������./P9v���đh����j�����
$B���i (��K�{B� �� �lT�"�����vHb���tS�iƠ\��\����GK���w*1�?�r%��_��Ѕ�O	Y{96�7m�K�hz*�O ��6�h��M9�C��r��%�[E�>�~�j��d�{�2u^��i����2�3�8�L�����xA�lC�[Wᚃ��N"n�ñ�b�0�
Mn������~a�I����g��� Q�߽����1�7�l
qu�3�]�^�_q��kNF��0T��l,��k|�eH�U�-��]��K�,�}l�2�O�l������-7u�n i0�x3����`�nц(���Ig����e����pd�G�0j܃���9\ȫ���Q��c�TM32"Қ)aR��L}��WX#6�i�FТ����Ch���2@��0�f������>��a�O�v4zpݤ�,��\�
q�t��ۉȱ/�&�27A���adf��n�}�a$)��(_g�ީ2 �aٓ	��5Vz���(�z����ĕ�$[��u�A_�35��+�H�t�]�}15��ӝ2���B��h�f�ú'�%�B��������� �
�W�5��o}N�)-qvh��|f�|��~Jr&��R��G�{����!%����m��3��,b&�zȼ��x6�9 �T����>,@��y=�
��m"��M����U��3L/�
)���#"���)f��H�!���ѯ�᳑�#n�Ñ��?��!���B�hP����B��V^k?�,�Z�_�C����PL��s@��L���0����D�q&�w��|^\#�.��T�q��nj���~�D��J &�f�l���d�i�������z�]2������y���dm+���򣮁h������U���AFuV�2�-��Ӱ�R���4�k�_?��H�or�@�S��r�3C�S��YC[M�r�����f��1����^m��錽�p���0�����`n:񊝁�7�pmRw� �TqS�����Vx{�박G���]]��O0����X�0H����]�n�;�3�)� ��8�*�85G�5Q1 /�;~ܰ'/ՈJ;��˭Nf�ɻ�!�J�&A��= v�B�\X��8����f�H�Z�U?�Y�a�9�<Gp�o@S(j�b�����0�c���D��͕	�����a�(f툮�9�����u~�;;���iF��Dn�D��V��c�G.uH*QF�z�]��)嫟�[����7>���ox-:`�bؓ��G����|`i}���5C���2�G'�܂����y?Ղy�̇,���o��V�a�����)1��*��IR�KF�s�|�~�\��j�}񥃎?/���?�a�nK�Μo?)�rFj�.���s�tbz�����q{O���B4�C�!R�x([M����P�A]`ѵ���ȬW�^vm�u�}7jO��:=��8[p�-�|�DP��`�R4M��x�����(P�������·!��\��Ч�����l+e�}6�?�.��,�S�+fN�]7q�P�̳O�������EZQ�>��V{���M.���ʋ�`�A�R�H9�
ďe/?G���w�'��Ơ4��{e��ō��/��&�M��� ��Bs�Ɛ\�MˮxBU��J���V�*�ԛq�ț�uB�!E�[��U��$Nǫ�Z�+���.mS��H���H��Q�C��X"�HD�M%]:�X�H��R��[+�c���-��2�\.921Z�1H�5	�nOA����t�Y��$���7^�&�Qsn�=be���M����d'�@7g+�,q2��5����L�8G��ٯ�"M���=�6>����YX��������4�\�2���Q�%��<ޗΌ��\I��������^CD�k\��D�?+rѴ�s�n-����hp�� ;z=ړlZ�D".��Q����Q����N�@.�#V�a,e�f������Y��v�v�p資�1�.���Ձ���:����T�n�w�yB�h}D��e?).h�����j�r\�O�$R}�U4�Z�������r���0�a�
�m�W��f��d���K��y#G<�sx�>#��ED"dx��79�������i�iN�|��=��mAc��,H�i�X�L$��t��:�H�V�j5��:C���7X%�� .��|�!���,ᕌp�?��&�i!� =�w��Of�RN������|��TC����11\1i-hܞG^9:S�M�����c ��ΰU�1��@�ކ�{2����B9o����z��������'���NG��������A�u-"��?�
���ɇU|�jH����8@�U�(*$��ȱn�7�5]�1�(�ᆁ��˄@/�c,��x<0� ���TWGVn��Z����j%�w��׾�v��D��es����/j�u�R�GD��s/;��/͛�u��]����`��2�iA�@�a�8؁ꐠ߆^�>���0�XK����H�@�rK�c���mՐz]��\���G��|��e�D�>��bϜ\}~���"��=�%J쬘Ӽ���|�;ԑ���v�%�wϱd~'�!A u��*��qV_/��v ����0�s��nm�������Rs��n]=ҶI>�އ"�B�ݱ�q��r�^�Q�f3+I2�{�0`�]���
�w�H���4����s�T�{��~��~am���H�^��.R}lu�@©U�~)-LG���4����s��o{���TMV�40�c�5#q�h���W�<PN���\��{~�)kV*ӆ%O�Օ@���.��b�<��e��`� ǘ" \�$����@���0�8�Z�&�}>~�$	>��DR+�+bx��crD�Qu��]C�`��'[���7t`��n*�<�Ft����H������i��|�%��#���5��CwwY�l�J�@�����ʆ�>��z��'K�ix��i�b�ī��&+$:��jKTAu�c�榓�~�C�A�6����f�*l���gKMl+��m���y1\���乮� ������js~]F@��s2�C�i	�n����!y�JAxZ$:!G�����K�fy��Rk	�^��"���p)�o:|cY�����K��e��KeG�Qc�׀A=�����|��Ȥ\���Wo��HJ�7���1>"X,Iۃ�i�a��	u��"r� �.{���224S��i�_jV/	3~7��4�Ri���k����6���&|���dD�y�Ͼ4��ʯ���s'�6H��&&��a����W�Z$Y�A�amd�rl�r��o�F�4�~�������S.�'W�r\����:i-E����K*�7�&�x��[^���x�&�|�Z臓��?!V��1lأ	����ZG8�LDVW�h�����-�2gQea�ZYˊ9�r"�.Q�� �������ʔ&��d��\㾖kH�����SgE����Q��Q/���}ۓ�a�E���Ǹ�Ǔm%���6�"�t�c�m����A-�}ꡈ�U֠�iv�0U����������>�E/X$d�px.���^x�>�bR{(�Yj�� �hx�bQc�zl�	>����N��0r���C��3ol���xa&I��_�E�jZ<��`��:�֗~I�)���Q���25�.�2I�lr�Zc���C�c��^ 6�ܸ��"`�EMx�̙�xW>���n��Vz�F|��r�t!�'�|U�;20�A��?E^%̶r�����cdF� |u�ű�����l5�ʦ�A���f�˞&���y�.G�_l�sp���a��=��?�G#���,ǈ���@:������ꭢv�i�2<�V��F��}7o��_�����E�c/p��5��C2Uof��iN���x��֬��(�q�72��1>6�[ۖ��~�8���L�3�����R�H�N
���J��iR�:=c��#�^T�u1n�c='&�Np��]Ҝ��_��i۶�j�9MV�>��ej8+�[z0�`�܏^�΄w�(�)���3���i���.!h���Krq 晲�7��"Y����`��!�U�h�l3�q��,!"�,��L�	�PUC�N���M����^���?�r�g;��Yݕm��i*S�1%�e�Z��c�X��`���&@�u�?��c�>��e �2�˄�zF;�]ݔB�J�`oҀ����]��j�q��NM���<$|[�C�V�Q�SVjD�+��MeK��x��)n.��R��A�K5�l&P�Tn��$AF�6R��]���kT�J%a�W�n�~��Rd�`�7��.*�B�<6O�V�-���8�)l"	��s��Y65㦏���dKM�,���[��$aw��z%Y��	צx�V޲�,�3W]X���k@6u��7������N{�����r+ObWl�o�U=sქ9태4<R�L�Զ2}�����:��w�)�:��ujjH�����'Wi|F�k��u����i.u��y�\��*갚�+ru���438��WLN©�K�VfV{��7��@S��a�^,�~���Ɂ���k؄�"/ő!"T<޶<��X%i[��X�5Zw7*��u��k�s�vZ���SR�8Z�L��Q2�?���Vt�ٖ�~p�s<�-�b:���W]�G&�Ƅk�s݂\u�w�2�W �C�p����?0$��aʎYYwf�V�>�S'c��Nu}J(�y�ߓ0�IO\�|EW����-�v�3�|�Xȃq���ێ$$�w�O�m1��Xp��SvLr�J��HW�2/X�U�T�̵G��� N������Bc� �m��'�>�Yx�U���>'��0�4n��M�Վ뾝��a�h	�e=�ekH2�z�1�Nm)����`�b֯>�rN�cv��@1���������χYb"H�?\9���[��T�F�Yج\��R��@.C�̝�q�� �*#����B�| �gH}�"��k����� '��'=G�{�Y�t���Ppډ|b�R�\ĤJ�Z���+�Yҩ5�)�X9,���K��TDD�B����������WAK����g��V[�V�y����9����>x��o�����K�I[�׻��O�F����I^��s�-�RN{���DZ#�a6�]�ۿWl�n�D$}���2���yR_&R��P���<<%�&���b4Q�6��������}��9��3��TA=!������?4X���2�UȠ?ڧ��VXrZ)�39��Uޜm��LҎ��h��7�B���A}�eOf;��*7��@&z��2�{	Ѡ?z믕�L<Up��bɯW�W��+-{kck]���7�O ���s�]y�`����*7��USSB�,ƴ��/&R����_���ܒ�I$����	˗![w3���aZ�Qչ�{��
P-�νdoh;�N�����(`��O��U��=\q@��ftKE�彝;��Q6j��횟#^[Z�����
�Xu͠r�Kܬ/���!����4�/\s��!�i�?�otT
���[�,�u'�˜����zYj�eDҤ]b���*N��'��sĎ_��f��$c�
HՍ�
?D���ݺ���|��~�y0g�ޮb�0��[EQ;�M����C
����S��W[�-���0��^���֙C4�߿0m�tn�S�ՠi��NBѪ�N�5�vW_I��-�����y	���se� )�R�-(ipB�:���ټ��,Ԥ1��d�d6	m0%	V]�X��@���Aw{���٠�5{q:0[O��L��E�̘���]�W�)&?��g�7
SMg-��`	 V:��8���=��g{ɵ�\���9<�Cx�ó}D!�������ͦP�_:��m{� 6OԳ�����?�VI�2a����Y���z����H�>s8{Q�rC/j���Hk��,����b���̓r~�+�,���n��_D��R2)������7�������`���I�^n�A�inƺ����xdQ�)��n�:���D�n���}g8ܮ�Ę����c��[VBm�kp�J,����j�Lj[t�2�W���}��4h"߻ �l��;�޹!u��aJ1	ƹ�ߢ�e"�w���X��i���$n-
�i逜��ħ:^��O+C���-yh�Z$�����t>Z�8�t�H�>��y�����o:Z��z����nu���ʒ�s3�w�q,ϫ.ӎ&���\��;�$bo�@!+�f?pv�#�ިV��Y��Dg����MT�7d�v�QƮ�f�F=�Rpw�S�|m�<r��C�����
�d��/t.�HR�G^gޑW��҉q���8D�᳈��Bu4O[�؀O�<���o�H�'�"���,M�/��hM� 
�ߒ�h�v�|M���ˊ�����i,��6H��#�.v�I�JES�*�;���'��,Tn�v�]):�F����<�#P�3U�ǎ"Y[�7i��Ս�}�!��ۿ�JI�2�$�[��v#j�4y�� U�gX�K�X4E9�VY-d��~lN�@���<ݲsRZD/]{=����iA���
���)���YY寗�k ��Th)I���dg#>������"��EX�4���EޙD\��m�.�������I�`+5*�N�Z���y��ZVwyE�8����xA�����3 q������9�8��f�PA�^y���Fr����V���E��\9�R����{l#;ZD�����^�T���zG�+~�`3��i�v^���@��zLtE<Zvǀ�m����9�;�}�q�p@���ﮞC�ȏm�T����:X�t�����3�K�;v��-?�c��,��.~7׺ �S����쾵���T�35Y�u@L���/�Y�䒂GK�sm�0��l���M��dbέ[Zq�{Q(����}�/�Ke�aN-I�(&h}�!�k{�R�?�Z�����Sq����"X�~#_�� �F��EwK�r�q���CIOʧAj�+&�k��G9�^G��L��0�B��ӕ����;7����)UK�C��X{�H�M;�=�ydw$ȍQ�FЋ�M*j�D�"On��������g��e�-���%y�j�Y�WCۖ�q�^	П&�7�Aٮ�#�ܑ�U"�h��M����o� c>�^2M��8��/ �
]���T5˨mf'��c M�fED���b��8������_��g�Ui�����(�e�*�>�Z"`�D����2P-�4d��&���B�CM���ʳ_U ��=
�"j����9�8I��P���k(߹O�ڜ��{o�������ȹ%ՙ8�֦��"l:�ޭ�0�޻[��/�,�hx�"�'b�
�wC��L|ٿβ.H�w����,���+�J�b;�f���:�E�� no��5j'��Ӡ��o��x���L"���땥�N��F�Đ�&�6K��L�!�c��9���`T�����B�[V�"�����R�,8�9��`?"|�>��a�01����C�ƭb�Q�"R�D8�ԕ�)Nu~�<
�_2�B b�)dx�u�}`jM��3����\(���i��P�ە��Yr���ޖjac�^��W��f� �5��R�Eg�CR�pi�G�	���ݕ�h�Y� Oa|g��
�6�.l&G����2�>lOy3��[���0��\\bz%�a����qhc���#g�f�:��&�����<�H틀e�~�t�C��Ze��N-��P�v���aX�����=�[PY�5��.��
E�$�l�
����د0��Tf��̝)4��:O�sD��%���	�`�C|�P����S��2;�����p�����$y�����}��U\��el�?x���C�� =���醣:��a;�7�'.��ǉ����v��6N*������y��=V}J�[���t���͞��1��O�C�� �󽝊A��P�W������G��I�e;��L���Իĉ�D��j�
�I�b7đ�G�����,�_����zF*�3����+�ã'�LL�$rM�ns\� ���cY��e��%�����a�b��Q��RD-�)���]
�*$��w�ǰ��X̿��c4N�,5F����8�6:_���8��t�o65ImvyH�,��4f�+�y4X���8�%)5���?���?x�~�]Ъ����""������s~r�J�0��wmJ���+WGL�a���H#թO��k4�i��Yp.�|�+`G\sQ�r�m��˾־d�@��pcs���iX��Xޘ�pʿQW�� $��5�S��K�8wfQ"��A?'�ȓ��iDR c�o�<0W-1��|<j�B
%�zܜf�c�&��}i�s:��$)��3�"��{�{GY�Q��v��~����J��<>�XEqH���''�	P8��Z���~���ey�X?�1�J_S��w9H�S�gu�����K�x۟��:�P��Q>2'����X��;H���a�9&�Y$.gi�&��~y4�g]���$�E�ۦP�������0ᡄY-�#F/%�aP@��,���w���Sf�����_C��d�=��@J���
ñ��Ug�Q�6�ͷ3W�ti���]�S�Ϟ�e3?y��O�4W�7�vlg=�ⷌ*9r����>�i�[�I��R�&��K�
~�Zt]�����nԟyr���!��
DE�h���N۞��|j~N4�et!�8k�Đ��ɭ_���� ����g���<��9����Ў4�h���l��0��{뱷}���̖.���J+���0 <��Xs�PC�dq�����-	�`FY_�o���9`�r�kY���Z�tv��+�wW�[��{�Tb|��n~���5��`K�KN��*�G^��� �`���%���mZCv8��<	���q��&�`O���#6?���l�ƙ��+`T��%�x�z�Ñӳ��[o'�~�$�gW ��:��.TÆ��i�V�nF���2U�p�RM7 �㍔QC�c���㶡��r�q�q:rG�c'Է*�^8x|>����58��&���t�P�o�x,#���}���
�1�v��t�ȩ��W�4�O�
��m9	A	�w�*h���R?�b�sjT���~�l4}C	��u����1����v���4��Q��#���r�	\��*�D�&�!��p��7�U�����|��C�޴��!&�V.���uT�G1O������ �]���.wMZpa����t���h+�=���	��@�r����x�u0w~|���� /�h>a�Bӧ{p�6��"��g�sCϢG��hM�:�#l��ǈ�fg\;lxi�R�z��U���I^����Q)4rWFy�H�OWB�Hc���~/Н��kNDf~g�1�ci�~��1��p���m�3v�#ȫ	^i=Sį ^ ^�
�H#V	|u?�'fm׫d�i?vbz�����j��4~�s`���Gq�!���\�֒�}ҹ�D�4$B����潜��L���7���X>�Y�y;��&*gX���H�B�]��=��asEY!��x�ך�p�[�D�ĕ�u�?6��$��~zqQ�ñ9&�%e��iK<pu`�6Պ38#��V��.E��e���#[���n�z�j����Z�E�I��-�x��=��Ǔ6��i��;���Hp�q�L���Ot�",ᕢٰp����G)����~4o�j�R�x*��AT�l�m�ˬzu����͉JL��[�|��^.y�\Kd�3�f<�:�#}v�M��o5t�/� |NW(�� �z,������ڰ k��!)쟭7��EH9ʀ�zch��:�ǵY<����}�1s]9@�������ҟ���=�\�'�K	a�R\��.��Q/6�!��X0�P�D�l���C�+F����A�c�ġ�[�����3ʞ{�?��-���̭{y����P���;Vqrr�>2x�_ ���%;��-��\�PjQ�Ӓ��iW�	�{�}z&�4��#�va�'z�Kp� �/�iS\RJ�Iq�C�U@$����.jP�&��T�dsrSK��~�*�,�Y�ϊ9���|�+�]�Q����nv"dV1a>7A:%{�_��K\W�	�&�(5S�<v!ǅ1�_�bdl�T���F����}V�/���~�q$Kj�%���'5!���[T��j������{\ĝz�)��%��u��Z�7��`1H��[�R3K"uϮn��Jw�W��v$�pꏄ���>�+��Z��UA�_���5ɟ5u��|D�d l�`�^�(i[z��Vw.L T�۳Z� M���?q���:�Ʒ�D��F�>0]ư.P�ź�k����X�-���T���|c�I�����`L{�ǔ��u]3�
�6��[�B%٦k��C��
4�-��o_�t���j�Y�������P۲'�R=��:�/�*�M��/8�B����M�
��3�Do�*�?R@ሱd4wf~I��1�s�]Y%���%W$ (�n�D>ls1�tk>��Ƈ�rV�0���n����� /����}�TX���B	��/n=�',8�`���	�}���>�"�YNₗ|��u���ˤ��:�:���B��y���B���#wm��s�PAٓ�"*��R׀yl^&T�(xg�w�װֈ��Y���H�^T#�\`|�l'yU m�лz�3C�a�V��j�H!�Y�������F�,<o�KDv�a����"�
��~>O����A];��wC�m�:����KGۼ\�S�E	$��q@�6��f˓ȲH�o��U�M���,Q׀��ί[Ig��J�*U���LӃ�1B��]��{YT�2*ȂO��<+���X�j�؝�;�b2���]ǀ����H�p��Y�@���"��=��Yj= *QkB���-��c��.���>���B���W���\� ɭ�c�W������S��v�Y]�9�.NJ�KX���K���K匛	D�g�ɨ���Y����?�:�W�*�;(sR���:���< �3�L��_ʿ<o,U�FO����`m줒��F�]���iP���7�&: ²�S�G��*תE�גSMy�=�62�q��ҡ�:HC $2@���]�m4��ܤ]�I����ᩂg���mc���d�=��`W�N2��!��?d�d�N/�{�Z��Z��Ӳ�S"|R\{ʛ��3�����(@s� �@p.ф��Z�@U4���ǻT�
փo7�w�����Ey�]��+e6(�����_��,���H�g�x�f�d���E`P�v���.z�4��$���e4�?�t�QD��dZ	_����]� �ȯ��7D�O)M�#
��)��H�p�\�L�E���?;���L�bQ`G(���5O�� ���4��o�&l��R_�����)q�վ��wn=�d0��m	��_��Ur�Xt�'v+�7//^�Eہ����L%$�,��c�2I쯚������|JƉ�!�7=5ZD�:�_��m��bŌ�����XY�8���p�a18/�L����<X_a!`-谜�
�E��!,�P��������k�Q�&9̢��q���G��$�%v(�pDו))'����HF8�s5=]���x���u��#�߸�M��{��~����`Vn��*�|kK,�����+�.0�$�CJ'\�ySW(�)F����"q�q���$�BHubZ����v=1� ��������& ��YBߦK����r��4���l��6��u�=05XnyB��Dv�R$F�k�Ky�D'9��^-�b�|/�z٤͘2������!Uu��PVs�*Hu.�p$[��� �	h:	���f�5����7Y��OC�|u�*̢�e��䵬imR��P� �9�B#��c�W�g4<�7�Kk˴n��.��-4,��?��p��S)F���l�UZу8ߏt"���8�� N�gj�	�z7���}��V��9R`�G����E6��2>�(��^��ï\���]|��'v#�X�v���x_ ��	�O�Ž�0Jk�+�%�Mv���Q���d�f�ύ��%U��I){��k�(����H'�Њ�:��6�Y�M�DE����4�o�1�\z��A���<�K��N��1_(�u0�$	�	X�jG��rf�ay�=SHi`,�{0O��AKy�c3�)�`ϧ���c9|�j��fL"�X��k��7���Ai���;C�7a��� ��3�l@�,����mV�"&8{�#v�g;� ���y�i>4����UM��9�[|0гKc�
)��'�tx��|b]��b�ߍ�ǲ�D��Z�N� I�IEp�De��撯�(%��Z;<:>{�mB�)��A查��'F�٬���A�9��8�icX�yz���d*Z�1�G�HBk�q�5���T��I�{������K��w:�@pD�: ��|!�����^���E1��LV!�^V	����zϘ�ɼ:|ڇ��$��py��������{wBtZ����<�GD����5��B-����WybyL90���:��*�ThH�)�M�#$��=LEm�X;�3�A˨u���뜨���!,+��?!-��_�����,WDX���8���)�����44�I�Dps�y��-*�:��'�PU�<�\���*����������;޷��|3����P$q�`���z� �n�6���?O�$��������U��� d�@������#�:����w�u:��ʩ�t?8+���5��\6�:ɉi�p�i*m�f��mIe��Sm,'��V-�TZ�U��FrΗP��bd��ĿC��a$�(�k4��6MY���$�d/-d��GmH Y��!u�l�!O�f��H�|��R�AEO.E܉�1T��'�$��;=i�����T]k{i���*<{-�/���$��ew[�k��xXK��cs�$;�E��6�$��xb ��6���5����݄}B��#�UK� ̢ ^�����w�l�i��|  x��7�@[��Z-�32�z�)�c����"�S����-�bvW*gJ[(r&��d#��q�̄Z+0��Q�)��:�wqen�C��������))�Pk���V�_���Q볞�c5R�-��{F^Ca���>��:��%D���t�	�4YK[%�l�a�����X�R��=��3�֜Μ�$;���ұǾk,b�����5ѩ������ץ�������i��=KIM��;�K	�ǅ6�#t���@��~)�S�,�d�z��,�Z�@;!u��
t{��廷�p#aKC�Y��]z�*�S��[�pMs[�Ĩ�M��6I9��~�Ս).��?���6�dl�|��޵W,���)!�5$?m>	���V2��M�S>�Po%��/$C���d �,��z�U��J�� �-ʶ9^�74��Q���y1�?��~(�Yi>��b�Y�� �n�M]�I"��g{>�Z�V���EWc*���_��kS�q������?j���_\ڇ�aAg�ox��@�C汾��4���f`+嚅)-/��x3Uc5nV1���`C��2���"�)�l���oR�" �����vu�P{�i8�֨R�R�zR�'-�O���>Np*ۧ��	 ,�[�|��%H�#�x����EI�j�n�4�f����?=��������mg�R�_?QZ��>��޸���5���դ�r����U'C�?��L,�J
��օ�a�T��f��%� t��-cЅ��	|��PnT=�h��q�^F���B����3�]��x��?w����c�[|��a���|�ܷa�����-���Ц7!�x�a�w[+IH{�SE���{ؾ����4�~�B�r�!��gems��A���Jk�r�Q�y��)|%�{.��-,�ꕘ7L%ؖ��(u���&��_�^�@��������|�� �e��&t��ַ�,���� 8D��;�����R������rx��%�S�bm�=ʷۯ=s#�����{%�;t�B��3�L�>�W����}Jr�'7"%W#O>��xyW�M'�����$����TZI.�*��t�i�������Y��c���}��2����	������0��ҢЈI��#`��8�6j�Y_!)�]�h��e4\��	��Gb@��~�
�f�������\��Qr"�幵�	����ZZ�&d�Ζ?}z�yrZ�[*f��b��&=6=ܖ�i�$�_��o^\�5+���&�F�+,�b�|��"D�D���|@���s�9�?��Ȝ��$X:�*LI�b�����#8R�mc��	��RU@���C���\�d��P��ecڐ��JԺ[�����v��S9�#�@z_��!��
��bɄ���|�&��k�3W�Kf,iv����	$��],�S��u�C����Y��}��;c��M��?����U���U�)&k�k7�m֠ŭ�C����`;�5wֵ��3a�Q��W������M���t/�ϭ5D*���8���@���d���:��y�YCP�a����D�C�L|ek� �ƭ�߳<��[�-)H
6)�>��G��|l�3��B�L��k�k�r�Z�ez�( R�=�o����R���`�fۘ3��;�]�Ì�&}���y0��qd�i�T2pg��0���}��b��-�v�@��,���GF�/ԸT�׌3��A?Z�]��r�Vꙸw5w�� 1��ݓ�%�׽w4)�9����t�� ~q�������J|ξS ��l��@�f��g��Hd5"�¼���o&ې�Ƭ��=���U�{�g-�g;9�@#�г�E%/��ЏD�{����o��
=4��M��1��qD;y�*���֫���d�;nt�0p��O�Pm��[�L�w`x����7�Q�v�X_T}+i���FW�5qĚ�t���_䘈LRڦ�Gӡ�́�,�&��Nn�g,%-�vyy�Q� 1���}�J�{,fY�~I�g)���B ���z��1$���e�ı�㨀��F���b�S<j�����2�� �$��=��taeD�N�D�?�����T�@k3�̤��ht��gF}{d���8?��"���c��Jܡ��ߌPf�����N���� {Zw]���v�K �O�6{�/�D3AGA�(B�`���κ�]I����y�iئ�k�%�謃5r#�Ζ8t/.-�Mtu���C;ĝi&7[��Ss����6��zQ@��[H͇�}<��{�(�o�9���/B��z2�ne-(����Iuo����|��IQ�`��i;b(��+Q�x�ڵ
�?��~ղ��ύ@����|]� ���jd>��*}׆��՗� ��!���SSg�/mNo���f�yr��x��8��o��*�{C�*�	k���74�U���Q�a��i3]'��aEȿѡ��������U��R~&��S�T���}b������@��� �Z5w��j�3&���c��z4�̬"��9�bm= צ�C;a��;Jk�Y�N�n��py���R��]y% �/�������Ը_|iH�@���ЦE�H<iO8L%	�^�|��������6#��e
���;�B�� ��q9��1g{�M1���-�s��%��7�]��f�mS�������_Ù]�g��)��Փ�EF������]tz����m�pW��醛���ˌ�GMRn�򘐽�x8�{BW�I�W��и�V�F���E��`�M�~�J�-��5������H7X��´�1�y��e�_L�g�����~�;m��4g�k�S�s,�}8ʻ��?�z��x�ԦAE$�� l����.=pN�G�dH�S��~�Ȱ
���>��UWBYt}lpP��,�Z����xI�>^x�"��CT���$�֞�|o�	�q̚K�P�!v/H}�c���XsB|r�a�Gn}t�`�����l�Щ�t�D�S ��_R��a�����������H�%B|0FZ,�����S������5�)έ+����mU$4��k� �Dq�)�=,����mй8���2p�h��5��ļ��
Y_��r]���xG�:Wb`�p�lK��(��t�h2H�+	�|$M^Ƚ���48f��ĒB/�����L��4M��1��10��|�ٗ�Q3���kte��e������^!`״�ٱ�0CG��g�j��@�g9p���E,X��.j㩖LPz�ۘ��>�H�5��|�h��"���L:o�xI{C卹��������8xg2o����-���	���K�d��J��xG��!��wm�J%b�
������ת�$;��ڳM������af&���ۇ:���ɭyg@��E.��P���C1�I�	N��a#'p2~ͺ	s�E�-�I��R��)ˇx�h��Ԟ��y�BX{!bidv<�>�*�=�$�R��o8쀷������5�v|�~���ֽ��j�T�d<�sdO�,�q�ve�c�A�D^Sthg�2�aD�"O[�=2J(��JS�i_�(���ۈ�}b^^�W�e3��"L��L)�?���z%Ϥӏ*o��:��m�-<u�iԚ�]+�K{�q��5�P­#��ǫ�W���n������UV���rH�L��1W�hB������]*�scI�G����R,2�����voH��F����:��x�nPr��J�������Z+�7�WX�]%LNDi�B�6����x�d�Q]��P����;�������gt��۽��y՟~��&`I���u�����t\>5|au�`"� ������4&˲Ԡ�y�`��x��� �U�
��a�a�>_Yi�* k�H�HQ�T�H�K���8��h*�T� MW��ZJ�~�q��t6�e�"�E� �ӕڰ9	4i�Q6jI��X+��Xt��^�>��ca�bv����J�M�h����7�K �8�O9R�Χ������� ���#�!�`����lr�X���N�:�a�o���q�f��Y�y���a��sj;�9��UU��u[1�;_4���P�p�zp�uT�j3I�Ui�:�F��Y��P��9�fu.��$.�WO��6,��N7`b�a�]�(����9�/�k᡾L˲��z��g"��c���)8�1��̈́��'&K£
�����	&Y����(1��~�,����t��*�t�د����~���ny4�����s�����<I���+4x�$蜐�c����%��.��u<�Z�\��4��f)	ҁ+{��& �F�Y�����-��%�^+��	_W�s,!m�Y�Ȃ�3`�h��l�b�Mj�WV�v��u����Q{�gڕ+�j��5�;K��C�����X�9�jn�������'������`6ƿ�o�bo}��rp�J+�d�"����ބ��a�a�|�#`0��C��=3�;�h�R�-~e��$�*�p��ʊK~��m�f݃�/.��
ٺ> �[�r�2�I��s�y�8��F���_��<
�)3KC3���'˵(Z[����u(�����l!��9���b���;��'��cU�5�]��9=C׾�#������V��j~d�Ȑ�<�v�IW�Cp��&�����ll�Q?X^,��w⾣)����g������Et��eȌ�D�3;bs�a8F�at0�7ƶ�[Ih�a?,LKI�3'Az�ȳ��Z��k�9G�h�b�m���[�F�|���B9�/��H�B����x1���Kӷ����N��۶����.� �����Ɂ-�i;9��3u�_���4����ۭ��K�YF��O�NpJ�#�R(�����^A�G�}Y0��
����kö�
-��]��Vk����Jd�5�F������3��v�ֵ+���,�Q�:m��gi�q��f�}!���cvu����F"l�	-
7$�D��ȴ]6Jq�Nj9:��u�V�����t�s��M�Qt��E�;�����б�8�g�M��6��L�E�~�N���E���w.�
�wRZ\b�z��.�>&�˖۹��̡@8+����
x�c��Y��>f��I�{'�����;TH��j��_�_
�V��\��U�	\���q=�)4i)����Ulq;�䗉��ohK�syp1*~	q�eڂ�)���ft����¡N�j��Z��O��|ܰ�p_�E-�¿;|�&d.Ey��";{��=��V|��w9�Jv6�j�3f��A�����?�2��: ZMBǛ��֝�5�	�}C�w�ՠ|��q�nȑSG��*�{����1:�N���΂N�_V8k݃	.x?S���]����0u�:Ɍ||��	꣣�;C�7<���j�}g8�����p.Zj���U�f�Q��9��LK:�0��	�o.�,�xt�/3�7NП�u����dT�И�	����s�Ryxw����lr�K(�|\����ў�	�6Qr�P��K)��m<6�fc|�bb�e%�
�}Ͳ0���㸸cЙ�2-�#��ˢjH���]�+\~ �	P<�>D^>�N*UYB�� ;lc�^�"�{��,�������j����U_,p�<�(��}��%��V�}h��{���Y|��fF�E�/��s}�-
p�EH���K�PQ�%Ց��,�~���E���y�h�-}���`�>S̘{����L��G�l�]���b�@�s9O�-"f	�q,c��\�����B]*Fc�*���>E���Mz�&���:,М�Q�^��^�[h&��ѴGB`��߻gD&���ά� m����y�`�\^W3S�O�UD[`���
g�tCJ�c-
Z���������1�9�z���~9��Xp�t����O�&�,�W3�kȉ�����^mp8��o42d�;Ҥ��:�ӶJ���'�M^3;������*KfBL��*� �D]^�y/��>vۦݱ�{QK������ѻ�Ξ����ZR��G��X�/������f&�>dj}q��{�C��fȀ�^��J������#�^�ǅ�rjLK��bPFaq����$�+E�2��x�> ��$��%؇�.J��)[֪����/0>� ���jg������{RUvB���፧�_[/�[� �M��M}�.r��w���ҋ�����)�%�P��lw+�pZ7K��;�d�]~=hE�n�x�]i��PB�&9NW��6;�!tx��L}���{n��i/b\�-D��?E�ēz�ʤ��PQ��QH��yv�L�������[0g��XB�I�b�T�(�Ff2q.pM����oa���k�\�A�ub�W��� x�o$d����C��B�rchדAk%��Y!M��	7�Z�+lmE��]m��35��U1WZ ��ĳ���N5j����ew�-�'�������U��҆�`U���b�e���,����ڐiz[���&���\�U]a���#���g#D}�=K�xt��m��976$�9�K��y���7j�XcZ�/�J��G!Yz��"�g�5��[-$X%+kGa�?&���"����RL|��N"����U��}|%f|i���顣����j,��Z��h���q*dM?�c*!�q��@��O���-XeB�	�/�7��~k�dAf�k��=\N(�Ar�[��V���g.�%W��JbqNY+	!KZ�}Ih8&`,��"&,}�Ā�M݈(�h�L�1^s�4�o�������Q�7(���L���4z0'����� L�`��¡F a�0��>�L���^k�H.��"E0��D2�Hxy�<`��xV=�{���M��}I��?��i��y.�����Զ���]�1�ᤞp��ab��M��
��Ct�c���5Kd����oSD��ql}O�����! �C���%��E_�=D�����P�PR��V�8{�)n�5p����^Wƒ\��4����(���Q���nR�|�o��M��R��:mmFS\�psK-�S����ga�M[ Y)��~Đne�>w�p�w F=����	K|���Y'Д��ni��1������7S<�Un�4���# RK�k������g�qr}���}�/O�o휴Z`;3S(R���~"�:F���{ύ%	v1�%����_�5�=y�9�[E��u~�����s��Y���~>ov�-��LKG��IZ��%6.��/��D~���\��Hɀ^�+�H�CD���}���>���l/��o�|9v�V�됊A�~\|�kO��U��GbB���tg�7�-S-	�.n���2��"8 �"��6�6��ΫZ9fmʕ��i�t�L!R����iV�9��#�/�˚�#Ͷ����[AxE}�@�/��)���̍�v��	��e{�Q��?���QHּ�j��ȕ	8��E'�҉���3�M�N�v�iz����<2I�L���K�~���Dr����c1��89%���oli��Y�0�:�Ҏ�U�:�v���z������>�T�a`пG&�����_P��RV��P��.����NşaAW�c|;���7X��\ޜZ/Vz=�)V���\V�+�ɒ�,�lP���Q{QF�
"�_��7����d�ƊIR=>�^�lWP#��j���;����� b;��Cs�=��/�M3V�U������N?J(�!�?�0q�6�óB����h�ڒQu���ޖX���#����p�Е���h�]��:N.o�[�`�l�z�[�y0q�?go*�q�O�����.7��39�M��O58_V���O;	�\.F��^t�#��a�Y&Ɉ|�94���X�,,
�&l��8靂܋����.c�wΰ�(7@��v�u8��i��X�kZ�:%�$^��2p��Τ��y}�ݛ�'�$&��]�%:�Ii"�\텼�Kˆ>��ҥ�@�"]��=��I�|�N_+�C�u�I .�����'�!�.�T�G~#�e��l���<98z��pz3p�p�HE�ΤbB�4_�(a07��Bcܰo˹��o��\��J���c�)Bp%ؕ�\��gY�!`_�����i&v>�M=��N�S�y���2��Ģjz���"�w�>:�> F���E�|�)��7��p����r���|a��s?|%ː(��̃&D�}b#/��C�;\��D�~ګOk15K]�s Hˌ��r7G��$陹�aG�]U�D���W��!��U��D{�W)��%�d��~�w��#�ϋՆ|�г'�kF��m��ּ���|LM��<�b�	Õ���%=)��hz�����)1�*:�m�m�ӪE{�G�-�է�����Ww�p��'�vWJ��pVfw�ND�JL��Ǐ@��pL���wF��ق�<���C���QhrxV��˵-- �s�\�S���C񁚐R��ע��6�5o����p,n�B\�i�q�oA%$`��]dr�&�&@����i:�oS�C��M��v��Qo�E/����u�w5�v�r��N5s^)�E��W�۸�����X:��3q5f%��S��'w�q9N�ٍ�-�S���i��A���%��l�Jz�]{Hʓ�BJ� fuH�{р�+�76/�����xU�㬝|���$�7%�E��P?�F���B�y��{=4�TA�!#|���E�h�h�O�Ç���)=��vBP��n���	����I�6��������lN����9�T�eu�#���w��f�d�ۖ����ɜ�X�{7����H`��B���/JP_��:O�cX(�މA�:n`��/����2�E,#�]��ʜe#S8b�rP�%j^����}`�r������C�t�A�[�+�kϲGa0�y�9!k��Rt��+�� S�~�z��)��8��ڃ�0l�u�;��='��Gku���騲�V���h�B
"����7�3g�=j5a$�;V����"g��śɑ�:���i_�gm�=��ۂ��_urC��3c֤���HH�u�R�kK֪��Hu������?�)[K�$�q�ɏk$[��q��SH�Z_r��CW��V�l��UK�e�����')��n�,B��'%|��_a������S>l�~:]ꊾ��P2Q��vaƢ�)p"N#�Y�y�7I�B@P�q`��<�4���J�0�a��yk+�h0�'��SE�]�j�XܖH�q*A-T�F���)�C8��(%:!t��g��9��	0��"�ɞ̅@�}���Ʃ��`�]��Z�< #[�\�v�hl�7�&����%���D!�6�lJ�h��PSi<��1���R�&-g��b(���DV��B�A.�J�&��m���w	R�OHv����9�4��ZJL��~�\<g�8�q�tz�P��&�xl���ђO�����T\A;r����LnW^�2��`Nb���J@��'�f,T�6�5��А�@ھ f�7+�������t���C
�UZ_��,�DZ��I�3
������ׂeh�Y� ��2#�d.W�}���jEn��	\c����CAq��dOuF7q�/k_k� :�I�^J9�yꛜt)l�F�����,��BhSPk9�C�힍S¼M��:^��M�2��L\�6a�<�z����S�k蓵T��Z��"W-�:�kiX&�)���}?v�IY�7��Ҟ�i�~�i����Y�;@�d�tvV7$�؈�$�ֺ2���F�X�(���� �.I�>
�:2L9�dG�艰�A�����@��0���H�^�g���h��/�t����CS���2�a,����ܕ�@���ړc>���=c�l�����4�{d�޴$����aH�A �f�G<�<�];�8^�U�Jj?�>2�xy��,�V	�pi��,�Ij��sB<k\ ��t��R0r��<�7����Dè��-�N��!��
�J+~�:(�_d�y���0_�R�vM�,+9kz��=Ѐt��p�\ȏ���ݞN&q@��A�3(����>7����h5'sx��6Ǘg���o�,n�ŋ���>�B�Uf��]O��!5��p�\�e�i�qV#%{�{���|f@��g��m�9v$&k�Y(����l$�݋R�LMj�Z&��J�Z��d8�Y����&CB\���#�؛�q'�l��9�;熢�����։�%��,�N�q������L��*yW`���kH�*/E�
�#�y�u��2R�JD#���В�H�ɟ�H�j�!�pY)�޳}-��7?�ʢ�J��E2��������x��[	u(����A5��7>��E��n�[�r�_�&���Tk�S�������C�#`���)����m'5/��`6ʟ�aZ�dA,T����҅�sx~�YE�N�x�!\�)�x;�0�>�P�ܪ��c�Ļ��%.�N��i}��Xsj�I ]rs��/�QV����O4�OSz��ua��S��v�X�S�~�Y���An�<��bTI �������v.4�����u���U�ň.qu�\h�L(�����Q- {\��Z��������X�l��<-�'�r��I�;WE,����ٟS�̸6j�$p�H�c\���\$�!R'���:��ӆ:cŔ�f���3)���U��h����N����r�-]g%X/3���-�W�8��G����ͱj�%v�1���{���3��E�����M�S7��'0h�篾.�[.�É��t9���kg7��0ԛ][G�P|pq9�;��8��͇��5�q��+���M�$����@A2�Y�W�Iy�Ɨ0u��+8������[�����M�AMD�Z�IY~i���#|7`���W�At��q����Y{�������|�:�ӎ2c����v� 1���x�	@��q+�����BR�� ���~�A��]~L��DvM��,���A�J24 ���|�P_۩XVS-��{��^�MP'-�g�@��4/C���coH4��y���Y��.��ߞ-7O}r��^
�e=� [T�����c�X{���ޑ07$"k��SЪ�1;C��
�I/O֣N��I�>�u0�.5ͱ�*q��]
{آ�t@�_8�,�
�aK��C-z�c�]�ޝ�U�Ǉע�>����ѳeŵ�TC� ��?���Ь-UΙ���&�~��RZK��mO"QC0�lby�䟷[7�B��%.���NX���KA��t�?���]sW���7�r�w��V���6���Ws���2IٓwC����5U���Θ�`����b��[��~��4�����r\v,e�J{�ڠх�3�t�C��~p{��p	�`��i~	�+��ͣE��:�Q[�Vȇ'��E�N�<.@�r�{���ϑ?*%g�&&YD�'}�Mbh�d-�Ŀ�~o�b�E::z�/=�� O���M�+}t%e/�s�>�@^��y�������]�Gt����Q� �V��P�D�������	�kFq�>&�TO�=�l�����eH�E�a´Xy[����?R�r�@e_Sx�n��f�Z�97���������o:LG��D��+��׽����R�S0���	�x����wk�g.	�MJ	d'�@���`�ЧYvbj�ÌzeV3�=��y�T��ӛI},��r�&����Vj|�x�G2�	�19w�bݲHYÕ����Q[��˾��nx�>>V�߆���+����?�r5e|tB\�a�6�4��h�~�ʇ3�8�����7!��I����L���N�k�CUt�E�%&�%�C �N~21�B�=bk��-d�)�jI@��N9(af:E��cţ����ͷ,��������v��W=����:�r�����{J�Т9�ɫ�)�A^�[���N�޲OJYb�G;ɲ��⅙Q���3�aD!�ܥ�t>E�{��s;'2�l���ڵ�'zMqN�4��j|Y�L�9ۈ׃ �N�E�di^o5�Ug��+�p�7��:�=��[����Z���7@v�حS�CG�&6~�/�D�u��>�c�^�IM���˙Ԛ����Z�i�7x;Ԋ�i�D��_Û2w�$0���.��#��tdb�py)K�(��~�,�kA�6��ם�������+��Pm>Þ�r��@�C�(�7�<����T;ߑo�J2�����&�f�������Y!�&�RfI�<�Γɏ�/��Rtp�5�?�%��ݥ�i{P�ܶ�>�xюh&���X���v"�l�ފ�1���M!��݋*��Az�<�~D}�N>U�NV���N�a��ߺʑ��%�u��'�m����A\�ч��P���1Oh�2�D��g���a�=0�K��\R���ia�Ϫ��MЖ�J!�����e�i��]Ԉ�+\�Ek�}p���M�cďqJ5H�eo���k�ս��5L��p4��r@�{:S����*4 �4��]|��`綔t����(:�B�r%z�w�s�O�2D��XH%�*^#�Ǎvi��4Y�&�)cź�����C���Y$��&j��ů�:?���JI0��m��"{r�Ǆ)&Eךn\F�줶6�4��Õ*�+~�/��+~�����x�<@\�V����6c��̚2�˭-@63��z�|ok�bdF��V�����o+G��K]���JD3�'e �I|��Eص�ي���~�:퓆 ^��%������j�����,@up��s>��/+ZO������==9G�����,1�h�,��lǄ ̎$>\5u�#X~�
��J��%Hϧ�f'H�܌������zS��D۠# \�M�I����'=>]�Ɣ�^iEQ�ō����;���S�3�	 q���~�c�	a�.ӹMVV='�D�eQ�}��Є��}�����͹	.[XYB��o�������>���\�]�1��H��A`�^�6E����I�3X�u�F|�� }ߕ0���t�\:l-���9]9g�����WB2��] ��@&m�5�pX��:��e�����u	m�`^ϯ'bdu=��Ĩ����vrVJ��gYL>8#<n���=w�2Ҝ��*a�Iu���N� ��	O���S	��I�n�S���[n�LTI�[�S���Hn�ƿ�u������?�fzB����Y���l���l(�}�0��ca�A��Rc@��t�	bU�W}�V~2�b�x%�!^J�q��mT��(r@U���*k|O��F�S�G.����$hW��`B�5�i���>�G�/�z���<��'r9��Y#-dn�@�b�$!��6r�|�=b��7��1�3���aT�JR��lI�:y���:��8�����,�A�qԆ}��CO)M1��t۸ܚ�}��.��n����w���tX�w��s� ����o��ꤋB\N��P���(,>�,չ���+��Y&rU�b��6�y�*����,9�3�u�},�]j-q�/�Vc���|���*e4���
�X��:�Qa#�Q���t]�o�GO���M�
)ge��Z�o�j��U�Sxܪuf\�0�z� 2���3,V3�Ky�?믠���B(���D㧮����q=���{�N'��hr�]*~o�r ��zuFO��Z�Dʆ��'=^�%��Ӂ|�Oi
g�cw�7Q;��aZ��V_��MA]�A�ϙ;��H_�M2EL(q��2 �|�@�G�d���Q�T����u���aB+%�E�a��Q�Z�� 
>���%{�Srd�P��Wb�g�(�d�lu�j�v�A�^ncW>����|0��j�-b'#��6&A��sIz8޺!�V�"R�=�
�>_M���`��b؃:�1%D[Xy^ף��8}�ÇC���<�s��Q�X	�3�ru��Vh(9�_�.�wѲ��l�6o����n�_�j)ؑu �lI�q�>��x��Ҵ�B����Zh�C-���<���N$�6p"g�{�	�hb��i��Y"�޽���CFQo|@3~�D����S�=}��ʀh?��ֹ�F����p!�=@��I'�^ȶ����vo#r�<`�Q�$eMd��]�)�gX�R�<����_�V���v��{�/;Ee �"������#nw|F���Q��E�Pa>!4�:���}�o�}�[[v��b�=�Z$�g� ����,�J�k�N���uɪ�E�k�e�#�	�<����v.x��{k�?1�+ex7�[R�F�W-5�e�8�ג��P����+���M��9[�\2Wt�2Hx�]�>=��Ư2^Z��%�py����V�Ic��t�7i�Bоvh�CĔ\ſ�%#����yj��
{V����צxǥ�-sC��.FHw��<1%�#�!�Y�Eޢ�jh�w�����^�-(�
`�����	|� :�����yr[	���O	�Ed EW��2���VԦ/C�n���W� 
 %�b�x*s�[��0�zQ
�א�VJ!�P���8��ɢ#6�	+4�ؿ�Xvنo����z���5[�Q0/2B��n"{�m
E��Vl*`OGB���؞�p�!��K��n�EU��FJ���O~
���na^qD�8n�8��V
���<��g�\@��)7(����t7<n��R�x\
�l��:H�
�Z�(q~0�^�]��`@�VLy´M���9����ĭ���ן]���Ŀ��cK-�-�Y��&�&��e�٠䫺�o��u^�ߠȿ��D����D�>icAy��Yĵ� ��j�}\��W��ݠ���g���������ʋo��c?P���']!�f��H�d��
���X���q��o(��k�&vBO=S.; ֭y(:�!��O�1#�;��QG5f�׭=1v��9m*1"�ȐOYh���w^�T��f�l�F�ȑ�ܣ�7E��Ťk�ѭ��F+d� c!�f�����i,	WͿ�7�D�S&�V�ù�@���(����$𿔷ֽ��	�sp�1���3��[xa��6�@�&�%k�	I�#Л���w��d��sB ���v߶�X|��NZ˺l�1�L4�snt��y�_��i��b�H���d_�:P�۾ɲ�/�n=��鮔��Ԁ\��v�oO�!�w�g�����"$zX�����t���BO̂ksW1̥2fJ��R~�,�|�/o�����:��N���F�־�%]��)�eӦx�߰
�t��EUT�)�U��|#.|0�X|�*t��L��.��g,@'N�Ԁ_�p!�R����<�.��KquA�JU�I��H�F�gcj��Q� 㣺�T$�p���Н��-i���t/%=g-��qo�n��Rv��/y�L�¿��h��;�0���Uun�+On�֒}��@�� ~��#CI��$C���HUc�eա:'%jG{y��ц�?�z��	XZz�&ik�0	 t) �\�v1�
�z:
g=8����4��tA��^�Ұ��`H��1h9>�RK�
'd�j<���ǷV<��+���k�ؽ����na�9��m33'��U�-p?\��-݇S9�lA�'CU͇ �Cm�<� ��4���e9�~ 9�."<��ZsD�����6ž�N���s�������s�xA�p��G�G-U�����J����{��yFa�լ����Qە�r7
��}�>v"à*��?�o4�����#T�� ��SR�������V+��ٖє�rT��&������ �IĈ1nSPk`�4��|Lw@(�o����\��eG�KY��d�).C��0���H���fP�hq�`k�w|�M�Wٻ��$�u� ����������K�,g �¿o ����5�&��gU��ew�Y���?���S�^��=n��j^e�/@�~j�K�T%���DɃ��]�{|��,L��XS�(k�%��AN���R��3���H��M�e"[��^�dM�2��:~o�_������[.��E�(�K�\J	A��g��ڬ �?2���!. �g�=�����0��~t�_�<���1u;���JE�j�p��k��{HT��ϩ�n8��9��d/�kw�l�.�����n;.'
��{XV_X@"��*���TQ��k����]!�o4�*(r�mC��k怣귿:=�q����	�b���J%���5f$XºW�2�&r�� �u׳Қ�K����[�d�-���[�I0X��m������=\~�}�c�s&D ��Ƒ.��{,e�+��t&���2�y�D��q��8d�2B��#��~����9�x�mۤ��F���%��V���{М�܄~��I�F�VI>�K�>?0��*��q��z�饄�"�P�,{z	��m�����Ef��ޞF���0�ݐ,��������9���p:Mj�L 13O��-���.�f���`֜�I�뭱��|&[�Â�X��OE˒�Ӏ��"�����՞�]Ҵcj�m�~vH���totG��e8R%]uy*��^�^A'ݩ�4��y��kb~�=+
b��`�V�'������#��T��Y�p�Q�G���Y ��NK��X*�w������L@C"&� ����VI���8g'Q���"rl���7�ʾoHǣ-5�|M��E�L���9W���q�?a凗k4�!�&��тb]"��C��[9jyut�3]'�8��|�P���X�<SA��!N��wZ������i����i'?-<և�:�'>���@l�5䌅��R,1/��	dkϞy��bX���-5ov�*��G�/�L������
��H��R�" � �ԢL"gN�R"m�2cn���*D ���_�P�nr�:�����B��{& J���-H�9#}V�!:���050�潝Q�~����D>��gG@��a?�Μ��臊��W�2�>�_��O+?{3�XF�Ƃq����{�NP	��+�:�I���s���p7�/O�v��g��=>�<^����`i7W�����:���� �M��H�1�&��!�]]A	֙���Z?U�Y�y��ޑ�.�7ĘO�C����g�F�z�&��e$��� ���]� ���i�����M�h.�k\�x��:^?d�ߜ��(ͫB���
���зWkSi���9y��]���G:��0��βy�GMp���OZA�&Ŀ0-�\o�kߐ�'���枂ؕ�� �SDJ诵u��=���UO�\��cs�(��ds씋�Dq�ݫ`��ўa��H���Zc�$�m�V��"ڪ2q�ſ��ā��x`;�4�X��6�~�ү(�߬R{������ʕUՌY�#'jm�o��!e_QQ��vU�i_��DN��)u���G�|ˎ�t�k��&�ۅ8(2P[֍��w��N��R�������q�ٮv��o��4�����ݣs쇠�����s��)��Ư�?v��q#��U�X��(�f "�.�7��Y�)	��[�,��>��#�31(P�K��Zf�����6��$�\+��o��P��J�Y)�9�/Ϲ0�q���WE<��5�B#\������|^���Z�a��w�hL�.ya�q�����˨�uFd�}66�:��p�����p7��!�ŝ���٤I,��­٩$���k�O妯�c��u:ۨ���m���m��P�^���]T�ﹰ���m�<Nׄ��`���R5"7�_��v2ȉ�;�<r���kg�52�`+(����{���`�@m��v.�K�)Ў����~���w7iKr����
�5
�åzm`5�C�>@�ް��;G\��}&��qȔ�3v�d.�4�'��۶�,�˯��c���[�����8��;|#�o���`9D�oR.�@Y4�4�#n���!��8�*��f͗�7PWh���gH1j�X�ۻk��D�mVVZ�V�"��G���!��k���L���K�(���'GO�{�=��n�ҋL�����&	��74C7@y�v�Q��l�U!̆�����8>M~!��\!b�׹M}�2������E��
�q�j�<�޸�zѶK�<-ӳ��"���)�W<i����� /�'��g��"z\Z�ԑ[���3G�d�+��.Ax�d&�t.:A<�u�\5&�X��BAW@=)c��7���!'] ����.�R�P= >&��as�,����&n1\y��a&����("�h]�fh���Í�Aˑ��,2A�Եٗ,��@/Z[p���3*��RP;����^}�:п��{�i�`��^�.gj�C]Zd�����ק�u��S0��g�OV�;��	�.������U7]*�G.��C�uw�B�!���Gf�_P�l!��h�.��n��+�d�Y�Ԝ�.��'0P�?:G_,�2�
[W}n�E���Z�,������)�8�'<x���H�4!ὅ�N�ñ��)h�sZ�2���T~f�/��L�Ч(��+��n׃y#����H�E���!�;Q	�d}������/�P����+#g=�XIDdU�e�o�w�?��W�.��;Y ���c&��	��]�����R�Hl��JI�[|���t����i�����c�D@�H��6�~���*b�����w#}sF��Z,8�J_j��VBgW?C�nt]������U��p�U�,Σ{n� �fŻ"�h���A�⓳����K]��F����JP���ƌ~��Ϩ(����t��%t�ry�v����~�
X�����_�O4��C5�A��V���c���hG��w��ol"�S�U��o�� ����� BN2c+$�r�->����NgX��|*f���0m�X��C-��
3��+N���}�V	�&�'M�jJ<<�>Ly��m�l �� &SP�31�]\Ҋ�/ �F��R��~��Kh�ɋ !�(�����ɭ�`݊~��b�200�q�����Nks��OѨs(6���=����X6�H�/^B���h~K�)��:��Q T�C� w�I�djFq./}��l��҃T���J�C3B�M�/b�0Y���� �SDz�K.���:���%�:]e��z4���W�42�&Ƣ�֑�W�o�J@�^���y8<V�N�4(�4̲��PM�͈~�E\S�D��Z�=ⱃ��6G�|X�0�����Z[b�gT��HA��<���>�d���$���L���׬.N ���(�
C���iC�X��7�����׻���[�w3��V&=����D\hHW=7*�h�����T{k��Z保�D�7��?//~p���)æ	��oAd6��Q�}�fH�\�:����P����<x.��,�(Ԑк#p��ئ�M��X<�݆^-8��G~�����@�0}3�n�;2\���$V뼒LE�F=[k�_a���h���Zѿ���e�' 0�3�:	��R�6�T0���c�Ԝg2�(���3��{�>ha�`y>凎n�l���e�it�(�#qN�o��DO�Nؕ�+��<���̡r?��"�X{�����Ǿ���h�֗��s�b�,#-�v9��}G�ِ�9��,e�	���U�P��<�'�̣�,�N�o�y?�%ܨ�^\�q{���8������K"��Oiz���n8��B��	MٴrD��:�U��|�,]��a`�_��c�"���)�Ȳ��N.QHzK���DF��;BxG^MM�ɳ�'��_|E漻�e�M��/,�P"��:�`κ�i|����kǃ�1e� ��}(�(��������#�7�t*G�f-_:m{�?��Aq0�H���#q�pZ�,\x9�Ȧ�������0+��ٶc�cn ����Υ���-� `�%
�ײ���sg=�p#g{����DFUK0��<o%}�L�o{��;�S<6$�\'��2�?��;��"�A��>�gx�
\���8m�!g�>R�*N@����uS9[8��*�4))0�#�\.����HN�h��B"�v:�$��CL<;@�璽Y�*45[�����d��F�>@�f=�;��H�2:W���P�~��Y_���%���RC<()�0�� 7_�^)dj�Ā��;�j����S�[��ZV@���D���y��ߝf{�ցM�k�ď����p],(bNe�o���&:6a`�OZ�Dz��v�N4�PH��>l�震�4T�cwq����6�t�y�!�h%�U��������̴yU�G�Z�"�\8��ҵ�{�@�Q�[�5�\E5-��f�LE��E�Ψ�P;�Y�����=W��t`5����;��>q��9����S��YL�!b`04f��nM���W�u�E��EE���Դ�2���N������cv�c�������v((W�K�!���(r��&`���k�bUX�b�ɚ��w�7�K��g4�-��Y��Q���7��Q !!��o{�����VǉST��q�%80�pUi-�dF�!����Ka8�k^��z]�B�C�"Hγ�3C�����R\;Kw`b:\��d��`Z9I�'�3�h�����̟���bim�)�+��b�3�p�!oYiy:��	Ź\w淓O'X�k�/��<yh���� ��QN�9�C���������h���Y"�d����$�a���o�u���0��Ȁ$����JOuD~�/ߋ�M�A%�5w! K5��,��찗8Lӵ�\/�c5@�g;M�����{C\1K��w��>�:�A�Ɵ��U%��T�
�	]�'�Jv�4��=�jAQ���	k�c�e��ڟ��l������o��.
e����g�D=�p/2"F����*��̤�o�8*y�ە���Y��;Z^'��!=���G��u3�J��/���G��.�� �3���dt�/�I�!��CR֙W�=6�:a�՚�-u�����8ao�ݾ�9MŎD`�ｅ}�Y��,�CPEd��֯�Ġc �AtU�	'��i�T�]V�[.��Ɖ���=,�ޜ[�iF{��fM3�2��j0���І��l�晣�&%�h:l5���d���/� �f$��V��s�$����@����q�͑��U����� �%�<Q��¿{է��+�1��][<�C��9��kKX�LS渓UVo0��֒�`hL��>(8�N`�Gr�G�7��ܶR`��|q������T�p(�`���Y�L˽��Ղ��4��f�e�~�XOޗ�
]4�-e?#ҲW�bM�x�[�,`��[�r�}G�X���ݾ
��Na�x�%�-al�
\��E~��%	Y!�$%�Z<K�i'��6Y���\,WK�-#A�XO��'��|wq�L�T��q��t�bR�S�=^�Qib���[U$�Q�q�궯��0fBWN^�����l�)�%�h-_��LA��W�vz��#\����ᕠ/}E^7r$�����I���"�Z FV����q�n�WrٟMZPO��F�훣��=�2B�۟��#� �	�
��	��aֳMb�����sv�%1�V�u$A�i�Z�jq�H�6~��N�5@'��]���dNXJ��m���xڣ,��б�������Ѵ"���>������m�d�+���RF?0���=g��S��?�#�a������<��В��K!��{���G����-�f����l�Ĩ	2�5�E_׋��tV�]���2�Q���0�IUT^�#��:*�x�rd�H;T��m{�T�Z�,)�*ʰ�D���8��B3�o�DO��N�4�y����rJT���g�{v5HJ�ƑU�s�x�%%l�����Q�/ОÝ�J20A�TAij��Ψ���xe�)*����
J*�$�F&W12���B��翯�Y�G��"ؙ�3.a��#-�Ѭ�t��g,��� 7o��M�N�"�d��-��V�3?�#���N�o;���?�˓4� #��O�
 �0�tz�a5��hZ5!�a��"�.�X���)�Ƈ�S���P�}�.���W̖	2T��pn������5��Y��%��8�A:��(Af>9�_tR������ˈ�-:�  ٕM����^�:p�͸�E��!�����[:5M�������I;���@�*MR�����z�*>��I֒8� �&,�ӄ�<�'Q��ZI�ʴT+��L�R����_D23�JXl�� �00Q�4{1�;���\�1>)t]�/�Ԗ�f�!��J|X��{?6i��{Xʶ�bЅ�
��xY��ouY��t�!;'�i���5
��I��چ`�v�^\�0uįh��(�~NJ��c�v��	�)`�%�z+�$��ݫK9�,�#ԌC.���:��ҷ:Y�)����	7����ϑ�b�f�y._[	�J�l�����钂c�gIItV�
���������C��xk�{�uv��7������hJG\Kj�1p�e��W.�x�v��M?ms��GaU%A���ۇ}�ם/~>
�`&�A���?q�?�����G8Γ�+q��:���"b?���G9W��F�$���=�򊬛[?��R>DI�^������X�ndx�����7���l%����
l���A`�!h'	�ܙ��]-�\�L�8(�֢���C���R��?H[!I��z��#�΄��:��bT2���TN�v����.�N@Qs��ů��Q�Q|_�1�٨�����ɭ`жh3�8(ɚ�-�	��C[э-i|������Ҡ��C��*!�L����h�N`� ��GkJH�C=��V'�G���~}?2��O��B����c���$�+�������oR��/�J���26p0������Q�ڵ�r�\��dE�j����=R�RG����bMB�T�'���k�����y�iF;T�������w� �{�Ĥ�Wh�3T�>��a�v%���ʂ���
!jd�kw�C(�y��9�?�T8<���M�uX��#{,Cg�m%�6�O?J�Y�3j�[��j���x��CW�C���1��vЛ�M��r?�u���	���彯{vJ�h�|{O����-�~;������PV��0S�FM6�����8=��9�+2���6^�A�33��@�VM	p���}�d�������FF<��W
��W�Љ`�|�ݟ�M�\#�i�Q�?��4&���Xs56���Y�{����K�,��S����CR_��0�4�1+~8�آ���d�g����*��X����m���{�I8'��i��9N~�qw1?�˯y��Y<k��!��2�h��w�sd�h��^܃腎0���.��
�t.�R+��k��I.Z���@,|��L��^J.�1z�s���{��H��5��[�3�Jy���_Z9pdX�O=�ҵJw:�z�R�O���1�u��͗-$��K$/v�Z�-�b�H�,�Ӟz�k��Q�.�#��	z.p��F{R��G�&@���TJ��E�@�L�q}WC��x�gA�ݻh��~yX2�I��U�zV9�00U&��B�/.�7O��-j��������4�xj��W��zꗯ�����S1Ge���S�3}��7����@�<�A��:��5�
+֗�5'B��4$�C��_z�w��L��+�`�d�|���£lC���j��^�puj�#0�\��?Z�[>�}��,�@)�tka�ӊ>����ؑVH��I� �$Ч��k�����=9V�rY��-Yģ�!^��QM�&��P^]�O�����y��zx$��c�K d�ۨI�'+���0�]�%�rD���^�\�]c�j�e�����d��)|�޽���T��D�bs0�&��UZb��=g�Q���12"b��c4��3g?�Na�� c�;
�p�"���;°��8�эܯ�PI����;����?��oN���y?B�i�E'2�A��v[_k��u����N��`���t�.uD��X�7qa�c�ZVC�T�lᤅ/�I@4��F�9g4�Q��D�.�a��?li���c�iS�,�s�1�J�px�ma�����>��S�Hu.��W��Γ{{��
4�4�k-�ݸ���JnZ���\�E�@�#�9
��|�a��"�D�\�R&��|c�b�r0�!�G�7������-w*7�Q z��y���걪�������ѓo����wr��Q>��q.�ŝ�n������W��jq3&�W��H?U���5�@%����	��:�so�����Z�g�&��K�nq��B���<s��ܓ=�^H��_~32��K�S�3�2�l�y]��
�8��D<A�[j �-Bu����_ �hԍEbg��N��XH��3<
S۸b�l����F�Z��U�F�0�YL)��:M)�J��:�s���<C�\� �XLZ��L�K��� 
�0C
�������j8��!H��G���Yɑ��]T�����!7e�؛_�`>��K�.�n�@X��݉�2���>c��yT�p`V>�u��S��F�ᔘ.�׮t��L�9n�9�|i�r�Ҟ*~�t&&��F����6�[aHv�1�!�O��篮��l� = �������I݇�#B��s�W����Eb{��讘c�3��?�\���=�s�	ww��҄K䲉�%����xD����N� �p��I�4�nA%������;�s=�o��yoo��P��kg���~�П��Y���`I�1=�� 3$�9�rh�g�0/%D-Nt��b��xVV����d���8/���=�Z��l��n,�;Bl��u蝲���r���N�ƴMU�����
^�*ᇺ��ר�֦����Mp+��Bp螔�B�j3_JGJ��&��fތ�aV݌��k�#��<v�����	���Ty=����w���fse;�
�[�#�drj�qQ���3��N�he;~!��E�$]�z~g�N�Ẏ�� ���}��Z��� *^���콳%\���AƟ�
J3蓫�ac�ʧ3z>�z������eY��3���"��=/ޏ5�G�$��D�ɡ�my�8�$�������W;\&����6��ۭ�����jYu��͸�M��/��s��wXR�L�Ȝ�ڍ5˓�e��g%��{lV,T5BxmT*�ſHq<���E,�V��l���bJ��:�}8A~6���k�����,ȏ�ð�Zpʌ������Q�ʫoF����D����� �$T�??���5���p��Ư��؄�I��Ɲ��U�v�r��z2�Ѣ�c ����	�~�[帜�g��EV�K�����J˒S��"��n4����,͢�eM!Ao#�� �j�p`B'�o���E��Q�鸀6��4�K��)Eg'���N�ì�aҮ��Sc�u�p�S C���b�;�:���}��uK'�S��:s:��J�p��_#�L^/��w��*��d������	���3��3��1�5�9K���I�:��?�y���I���0O�$�V��I���u�VB(8��I�7zh�o�T]"(�)�.{ܪj�Is`|��R4b�ס��m&y�[����u�}sZB���
q�	�gDݞ�X���X私� ��0~��W�VJ�/����p;%�,Զ/�V9���(�X@�NA�Ɖd�`e��?M\4n�mg��|�}��aJ jݍ'���B���VB$3��V�+�v����Cv�F0����܎�2�!��~�.'�K�+G]Ǳܔ�%�-���P'P��y*KX����rrMNe���:4��UeIw��	=�"j	�u����O0��b�����@+���>uP��b��H z�����DS���4�ͣ�m�^��ˡ�fs�^LIV"q5��#�����Q���
nG|L�����c�$7BO4i?*P��d;ɳa�SE�ܽu�����.�$j�X��Ҡ�'P_3��%���D*;��U7@Z3w������~���)�ڃ�F[�k��C��B�>Z/{u�����Tc� ���A�թp{��+��6SL�\�#�ر���?��5�7+U��K���������L����PHj�ʗ�]7�P�س�"��f}%u��J�N9۞�<VI��k<Qu���j۪�m�x����;�D�Ch�¦Kq���7@H��_��:���گ�_��,������݅���������n�]lõ� �<ff�EG:q��HJn�KL�����|�e^ǿ�d�$&�����f���-��=e�8�M˱���H��~��hQ�Bo���Bz&�]�@�k@�E+��>d��=�m�	7X^G�4�eB�".:f�AtZVv��k��x�O��w��=L��j�(�f��Ghy��0���{Sf ����F���)��4�`��k_�S}P=�S��U��ժ)w�JfO�X�����&�������eVt������{/g��7G\��C�:!�䍡�L����v�W�eP����]��"N0�<*ȣ5[��Ut�l6�O*�	�cDC{���1���3�cA��	�,�|a����H:
?�������)��邤�a&�q�Aw�_l��������+�����h�ϕ�R=E;��Vx=�ѱ��|m"�}7��Q������C�DoF�&#yC�������j�8f,�oi��7��p���)����/�APofƬ�����(ET��=ۏM�M�y��HI�vÓt�ѻa@�J5�{�%6�~W ��a�_yC���I��.�(�V�=#h��9C�S��oC!�4aKM���X���U��S���5K���2Vo�dص)/��>~����õ�����5��(N�	�MN���x��&���ԫܱe\�_�"l�u����D^?�U� ?b�ɀ̽x���_�Ii-@���xV1&/B�b�d��!���.���M	�[�r�nnu�i�4&]͠��z�3��K�OX�$ўw�~�WS����,M}�G��]v$�u?�լƷU.���dW��,�>u捕 ��r&+�T�]N����˳� �vtN># S�Fj�3)H�b������ݝd�g������s��#5��cl^vQ3}�3	���4�S8NЉ�yBo��\ȶ$j��tO&�O,(�p��S��Q�wQIBI��ߓ��/���f�p���(��n7���7m�g�y�n�0�;9~�G,���`�����H��nD̈O���跤5���qz�6sX̞�V?@y.��:��J5��S�A�4�FR���$��	��!��Pz�V�����V���c������b$�&�p�$A2 Rڭ����?�\�Q�L�_m}�p��!m���x�?��7o֙�-m�<�bR���F
մ
z G��Y�!��-��"�D/��I�3��b��X��W�;���C�8�(��Z��FNW&�4�*����p��t���%Q�Tڮʖ-�SI�.͙�)�e�%5/w6�9�R�Ach���[ltV������;����wC��]I��Yb�V?��#P
|Ɏ��Rk�ٵ��r9M^�`G����~��Q�@�u��0^�Պ'��%����t'���X)K(y�[~�=�H�x�	wR���
��Ξ��j>f�~��߷d���$M����a0��D점~�@� e��
�Fo4J����zʪ]ϯ��g0�3�+�j)����{%h���

x��J8���Qt���0-�n)�I@aV��y�8�����8=[�:h/���+���Nt���������#������0�}/�@�<k���ho��fF�����:M�������J�۸����3]�]�4HP]=���@��VaCr���-_�gx�-�q�]���GȚ@�l�ַ��Ĕ��,�h���(x����y�H��u5�-<�|����G��a��S�jIʮ�
ۖz��伧5��w�_�+�m7*�ی��LI��'Sħ
��k��2�K��E7�-䅒Z�=y���V[t��5��[0_QkcJ�gIcy�J��o�4���RSčjt��_*�ii�I����1$�z����%3�i�\���ȟ�i���J���ȋ�Ȃ�����f�S����#�J �k���8GQ�P�����?�E�R!��[��R:Jt+���:���^��6��ɐK�
�}_u�8�hn׽���~�'8����*�h�<�ΑV^jMu������_55A�Xb���T�X1�_����y8^��%�A�RΒ�ԳրU{��Ӥ��h*��TʇO�z��\ ��XI��-�|���s:G@����5�^]���38{�w��8�B����~�ʘ��hX�'�7�����=�/3�����/_�,�>J��
�����E�U�쮋x�Z�X��f�4�y�`~�iB=и��ݠYwS3(3�B.3�x!56/��Y-EB��rx�F��:ßP��"F1�~��U�"K�Ø6r��R�#ѳB���Bbu�Q�3�r��R�k�GD��n�k躀�)B5�DeD(>�F�I�M�h�c?e�>q��h�زȾ�G�<Ț�IYa�1�0�)��]D�& �r�B��9��(f,���ٞ�˪Z\��z���qz�թ��(&T���@��0%���F��	�g��4K�QpW;%�13=G��`�$��-�V�Gٽ'7 0A7�e%}؜���,;�\�ɉ�"���)�1��,/u=B^�R,�ƻ)9ғ��Lj@T�3$eE���?G�3�����=b&
��ncp�2�����*:|$��`o�W���� 51Mן���Q���,X�n5Th�)C�C�P}*'�@����Ko,�l.41N�c�h��j����R��� ��������<��� �!(��*(-�AR�KW�����V���b>h�&)58��i��h���F"v��Ӽ�����0�@Z^��m~O�f�q >Z\�*Y�gͷ�j��g��lz�CJ#���$��_N�=[/VQ������AXfd�쥂"�M<�����-� ���ӳۑ6�]{WCDG���ᐕb�����@�0�'g�A���-��B:Y".���s���__Rӧ�[Uf�A5Uɜ�Ϙ���JԨ�|�t3BQ�ߪ�S�{*���y	5�m�Ѳ�N�ÿP��^ϯ�DY`:���X#�����2�� �<:,Ӭ�ep�K$��`pCKHI<�J�Sq��,�����cr&r��\�(���_�J�4�p]Qc��yP
;�K�V��F�AК���9�җ��1�j�B��=�)���9.��?�>�3w����'��X��,�Cɒa�3�+rjK�	t�G2�&��@B�}۠kaK��	��pc&�f"��e�wd�ѿ����_z!��zGQ��h�D�� ��Ob��<�0��uY)�$4���R%�|����!~���m�"���&�,��'A���l4hBp���>�3�J�J��rqX�R��}����"���:���FǺ-2�)]�!u����G������&�*��r���9U3����L�b���S�
v�J����??{��h��=Ur͚M��,�� �Q߶"1��r��h,�!Y����ux�:U�֑[
� bsDl�"�}�_$��e�����bM��vp��Ck�ڍ�;��ixX���m�H��'�a\�ּώ��V� �mJ�Kl��8��䕠���fҩ�0&`�Q��/�V|�i�"��7?{Z�	���50~wU��C�U�X��<���ń:�<U��� .B�ˌY�0�)F���������C���g�'6�'✛�����y�P����2�۾v�L�%�^�)	$�% �_D��:�e@���ֳ%�x���d_���p_6Y�ϺpWE�kV���nh���h� ���φ��m����8Z�s���N Ҽ14y�,p�{���$A#CSؾyy����a�fq���z#��p2��/�>�G�X[����nG~c�=gW�b5\7�=��_pa�����g��j���_����k��n�/:�	����DuO&��V��_�	��8���D�I����ܑY���m�i�;5K����|���1�Y�s�|�Xfgɐ�Q:�W�M����ȰZO@���@&ا��;w
��?b& ��~���h�~�HH���b�^ Uǡ��UZ��am��r,5��u�{=�9P����4l#�˂ �HE_�{B��+B��p�P�_�A�O]��O��[*�7>�O"jC{�Tn	,�_ �Fa`����B�0 �kd⃯da��|�fi�Qc�݁�)-����
PNQ���ަ�S�hG�d�"�JHP5@�g�|� ��eYv�%zeH1�C�/������ě���ѻ')����@����;��HF7�
�}�	{9لa���P�*������hg���o�^�
T��{�ǂ,�T�j���<ihɋ�?uq���F�;ՙ���� �E��,)��$�m��O�P�:���ȦZ� *zd�+.���4_�V��D�NEw���ʄa�A���f�F-��P����pl؏]>вd�����\uO����)v�ǂ �Bn�#�K�U��]7�EW?�6�e	���AX��h^a���W� Ǉxur��}.�v_My�(f0�9-�������*I�5�W����E>-C�l�[}�U�*��Q��W�y8@j��pr�GK�!�.�%)s4�GT�/��!��;X�j¦@��B�g �KNݳ��p���x���Z��d?j�Rs�V%�u#��|B/%Z��7��X���p�RAw�t�8���$He���YT���4��{�]��.|N��v��s ��*ʞM5��9#OJ2�TߴR���:��٫r��s7���M~�{n��!3��wڻ�d_ݟ@�M_��K�{
�5�C�y\t�jD�i)m4���@Ҝ\|UR��񁏀v�q�:�yvbζiP3�b�|�[J��thKw��
&Z�F׬Q���U�R�ێ_N�@w�Y�G��Z�y���w��5��e{����GG���~��[�����ׂ��� ���KSa^H}hi*�I��I9et�@B�"������B	SS)*Ѓ��߃�v��Z,�q� �O�66��F-��ڧ^4�8L�W+�l���t�1�;��L����І4h���Z;�թ�.�����Y�N<H���n�/����{E�X w����*]�@� g�*dzo!s����]�B`�)�r�s�E��-'��)�1�֬�!@����~w�o��9��6�8�5×d�����[Q�}b׍�"������ur��n�.��x"�D����Շ��0>�ќ��e�R]�.F���nN5�+�.e)�����|k!|h�*e�J����
�Rc���;9yf�-�!ڲB����MGp�!�'�3D�����n�F��ǳ�����E Y����t�����9bm)�����4$}���12���������a����$fNMà�X�"�RyB�}u���65:�����<��4�F�Q�����w�l���ƪ3�x7����u|�� ��g=������y��W��U���^]V���#p��-��{��T������z=�nqK�&Bc��W�2��`{Ha�Ժn_��WZ^����>zP1<����|���l ��2xz;.i�MFY�Y���0Px�W��d#�g�tװ��{f�H�%�Q�ݤ�`8�������h��֐�� aۧ�|�R�Ӵ�9�YEo�@��ƀ���OJz���5u��n8 3�+�[�@wʘ�(�RS�m���[�H����^\Ǵ#`���e���⥫����
"ՠ	��EJ�V�J�/|]ݗauu@c��*��cEt�y)�b����8��Cu`X��$V
,|����j��jK��l��X��y`�,k�� A4N? 8�zדǡw��e�ˡl�����HF<+��D�}r@�x���{��$
�kl�g��-WSF�J������ά�ri;�z��q�wC��EE�b��"�A1a��
�S�lX���#��X�V��n`�%�n���-�j��d�:6j�V�Һ[����,1��3�Rþu�G�*�ܬRE�`�{h}aZ�X	H��
��kEq�����Sz�S�Y0(�I^xc��.�"~g�&7���u�}Rc���K��Zcy��Gu�GG���Idt�Ә�.)��)8�w7��~!��z���Jv,�#�g��{����N5v�Z����^��R��u�a2 �^0,��u�Z\Ӈ��Հ|���h�~�O�@��d"fL��}���%E�yq%|�s��]>��0���ό��eU��;�\�.�^@��r~+vb��2T�G�@f�����:	{��g��v?L�:Yz��e�S y����,V��W����f����P�
��[������XҬ�nEJ���w��y��b�ug�b_Cc-��pH�)�hŸ��(z���Wg�X�ȉ�����am����qs�g#��@@�?�AIĐ�kj��j��8~"��`�dg\K4�lrd�OO�Y��4S)L�?���S�KA��|j(Ѕ� z�nϴ�>���c���z'؁�Hk6T�����~����w�t�5���~�X�	T��߄m���dtY,t�4T��f;��$ps��R����cM�~����;���M��L3��X��2�����@�=�ᮺ�Lqd�~��F����,iT�<O�����w �y.��CN����V��ȐZ���4,���_�"�jP�uf���l:hj��_�a�3����ו]�S=�F�{���	&�͖��}L��^>|��+c;��(�DƼ�8a�o�+�!Xq���mb��� � R:�y�S�����y��>\A̪x�ijL9���[�f�˚���_V���ET���&��#�gS�ݒw��d�ۈ�)��w�P��i.s���u!���c�yɍ�1��\NÇ�E˝�/��Ě����ۊ�ݼ�<D�G\$>�S�~|���+I��?�]	�@��e����9i�����;�u��C}(s�M�_�4u{,?V�{y� 덟��Ë��ݵ%�- �b������b���H�ⵋ��u��U��gB����,�6<���F�$ؐ�_�UK�F�e��|8�G�^,�
�[��)T]C�?J*>Xv�)���FAv�4�����!��,X89��F�'�b2�4�
��\��qO�a��R�	A>G����M�6X��.�Ͱ�#s�I�g=���F���>�Aj�Q�s
^�{�a�[�
��1��ĝg�P_�M\=�1��x?V���%�߁�Qِ}S[%���l{7�L�iQ!�e$"^�Ki���K]�i���
�Æ��k>����ٳ�J��*�И���%^��Yf��o�$����&�S'���\t���֊NtJX�	�I���$�~w�*жf���T���ap/���W?���O25�~a�3>���S��O����N��RC	�I�ꟴ$3����+u����Ŵc�ǻd[�G*#�*1U�~bŨ�ާ��>�J�%ե*�]��<�^�RL��	�t@����u��.��5��d��td� ۂ�۵ُ�y8���&9�Jp����x�3n��w:[�nʪoJ���+`nlRmR�
�����LX�Z����s�r�l���D�=7���X�w�>�?J��8��f�	~^9(�,��Zf�-l`��؞賌Q�G�D݅;�=��ۜT5�)rY�<�'Ran�c����>�w2��ƴ��{DE�N��'证�M�����>���z�",����r�Zړ��y�'<����L�Cǻ#�J(+,Y��rWo��P�hp:
� #���^]Z����/����8�\'�V�T�8���d�M��1�9m�>?��2-t��,�*6���r�>QH� �9s��d�����lE �3"���G�cD�F{	�;b
�mXv5+	�E�Kk{�m�\��F�|��-�F߀i����qTx �\�U��X3��чo����S!�~z�]������#׸��0�gދ���B[<���GSU5�IeF��{U�RS��i%�g�]��!q��ʔҗ�<���(�����Jw%k���b;�����=ėd����Ra�1L:�D"�Z!q��1V���anB�+��k�ɯ^P��������<8�y_��~gD�N�XIp�C�]�@Ų�CM �x�C���������ٿu��*.ö���	iD�D��R�,�������NZ;-Aq'Ԩ�7V-`�s�}����!�'�K@�r�AP }7a���CU�V9ٱ�el�m�V2�|�:e;N��Hsw����p1�^ц��\2(E�>J�,O�ֈ���>�d?���	�Z���t��B��3mx�G���R�WDI���t"��!�a�2��iz�&;���
�ݧ�r� ��;�E���*����'�I�~
�cFͲ���`�]���F�e �q�g�Iu|(^ tH:X&�(��ї�$����ꭄ��ka����-)l&x�h�#D?R�<��\sWo�Є|M���N:�H��v��_�\hN0�ɅX�I��S�h�������9�����,!����y�:A����C,�_����B��g�}�ˌxu��_�]�_��1�.@�E8��ѻ�w�� b -����՗Q�����AJ)�V�X0�+�z���Yv�7V�F�*=O����[]�b��)ʍ�1�a�ֺֆ��K�|�Ɵ�q�#����0X��	`�����S)	���O4/���Mr�����#�0CF�*e@#��h��:F�����Frv疚br�r�goͥ��nG�O��5L8x;�9��9�y+�P��"�L�҆haGYf���"�NX�'R�J� ������"��pcB�4�Y%M�́�h�q �p�%�Np��8�sc}����ޅ���*��_Fsd�W~�߂4n��]�����i��͏ǵ�d��Dn�$��wH- ���T�]�A1�c(���l)��Qܣ��H,2U�G+a�Ve�v]H�b�Y�����½ ��:�z�=�O�q�T�\ݦԛ�������m�H�64�qA����:�-e)p��ސ���],���2[^UT�Y�g��P�Y�*���*8(��;(^s������yG,+� 3A����� ���o03'�&�Nzty�2]�����{s@P_g$��h���}~�j��8�ě�ڪ'�BtN��<�)�;M��I��Ǧ�)y�z
�p�"q{Z�[b��5JG�{VL���*�[@L���+�IXB�k�̰tT�3i5*@N?��h�nZ����$>��c�vyb#C�Bƙ׽���V��-�_���ǐQa)�9�7ͬ������f��9����H����� ���Y�:�LN��`��=��5��#{�6_0�ޕ��7�7����w���(��fL+�A�L9��ݎ��:��+�U�Q��8QMnǉ?]�n�q`�$PI��v�˸�b�(Tʾ��X_F󒑉������	�X�t�*�����]XS�^eQ8tU����ڢ$��G��]���x �z:��ؚfT6���O(�N�.7����]�:|�usxޡ��ۗ��5O�_N�9�."�}o�y�<�I���_0?��Ǣ�s��b��B������^�8��ǩ8���r�8g��~m: ��=hoW��D����y[�^7�W8[0KH�?4Q!lT�sI��
׊�|a�a��r��d	T�A��#Z��Y��4Pd�gW�v�:[�ɇ���a�7�Av�4gՔ�y3'����u������sT������0���Q��t&�.a�k�� �}*g9����~e슰)\Odб�tM��U����t��\�$o%q}}��7����4y+���/`�h#�,�T[g���sj����(T�C�żp��L�e�̔��"����Nɹ�O`��4H{�E%I����YxĘ�`��x���iV���}y�q2M�N�J)�P�z������5����e�s�ȯ����s@-63*��*��{��+u���C��i.�5�h��g%�@/���6,o���y�a<�*|ag�M�ZCb�s��-����땞����VȗY�+h�hE�+%���TMI8��I�
�*�����O�߲�=�XJ}u�͢���m��������.|}s݁[�,�����9l��_�N�Oa�#�m�Z�'�����~��ecW�o�3�&��:��v�w�Lc=5�'VR��R�E�φ.V0�{H��]�gT���(�����O�(� _H�x�w��w&]p��3C_�Y����n��6�ȁ���E����L-�C`]��E,2[3z�A���u�H��q�X��z3��V�ƚ� ��"���^�-z҆�J���֙7�{��P�t��6�-9A��.JDI��(�"���G �#L�)�.���i�~)P�҇�=��
�8�����=lY؊͸��Lѷ��4ȥZ{���7mC����.5p��jr��-�/�C6i�6��}��`��֤0��3Z�Y9�G�Z�L�n &�k�6m�~�Vv��W���[�pZ���f$��.��`��#:�S?�u=A]�6�)����f�'�������X*�a3L�ĉ��w���K�#G�C�/�8�5� !
Tr>��� ��9�.y��ky�e��=~RJe�$�H9�]�t)fT�Y ��(�}��P�F�Of��&E����?2@~�X��+�����"�#���;�����~��f�:�����
�@$Л��VB�I�Z�^����Q�_��V����
��KQ� �����(��	��<|P�g���Ɗ�2��y��	� U�s��'��*�$,!Ag
]YsU	��0q�;s��HY�#-���(��s��:���b��g0�L�L�G�'
/��� f��>�^Ap����M�����ٲ��OϭR�X@o�������:*(��[���#N4�|C�}#E]�&D;AP�!3��ˏ�V;�i�]��'`z�Y��+��2T�S[�����1.����CmPR�������@:m���Hw���Y<H���%����O��}<$:���P�i	jzS���UАY����n��G�CfJ�rA��;k��ک��b�D�S��[���,��RC���&&�5��"��ID� �Z��/���������S�)|`*�?i6��煆��8��[�s�����r�`����P�3r0��Xp\����i��'��\�������F������<��\3~�~��V;�n�*�1s��Ǘ9h������&�rd��D<�x����"m��2��Q���l���C��fճ���pq�f��.(�r�)���
T5q���ʟsu�a۶�Ú����~��폤�f\!����YR�J����PQ��ޓ���w��Y�����5DM�0���[��:������ ����~
��'����㓉�~ ~g,��o���G�_�.���껴�"</�\��1��e��0<�^�)�$Q����6N��4Frxź��lNU$�HB��KT&�݊W��N��k�א����>V���/����N�d���2g�òg-�ɜ�g�j��~�MyL8z��H�[@�ٸy[��V���}I;��Gg"BV�Ḙ�����0��Qi���� r��̰� d�xx��&xn�z����F���~�^}=���v��71r�:CDp�ӗ�F���N>L��eh�<��6)2fN��(��WRuڹ���2�,��+ �%�_���Z��E�d����#��V��]����r㔩/W�;�34�^�rV��o=�}�k0n6<={����	�릗��0ē�|ۀ�X�2�5R���N? ��2~¿��u"_��JG~�4)��_�v2���}b�����Yf}�o��>hR���H�2�<�MDx8�~�C�OG�$��q��c�������`�&�K�U�X�393U�i�Ee:}�pP�������JRr~>!�����JO!��q���F!�e�#��f�oA5��0�53�$O')qT+pn�0uH��k��{�i����	�#�Z�yG��񋾛��|�9X�M�~	z��k}O��V�;�p��y��	閗��5S����d7���wa��[�W2��juä�fi��G̚�{����i�������N�2�����������fs��p������n�4w`M���W�}�g��!lOy⟑6պRL��͉S�����ѿ/�B�Z��CTz�e��<��fQU(q��px�j�rzV<���R�}�W��4�#�d(�i��uQ@�a�]��q��"`�ꀍL�_���|T;�.k.��|8�F�]�婱g�k�v>m��ɔ��Ä��R�(z�-�5u�®/��h}/W��I�Xߊ߅�ݣ����%�@ޢ6���%o����8��r�f�}(�F?��� ��6E�����X�`oP1v���y�ۃJ��;�������(*	,���x��8���5���V�h$��tf�����+�v����x�}��
�M6v�����W��Oi,���:I�>�4=n��{���Ǟ�7�f�����T�1��	A K�[�.��A�f�� Qo�f�^>�E����&/?rј*�~�z!uō�2(6�X��	G��Ս��=�7���w��@�D,��;��KC��� ��P��$���숾���?!(��ݢ�낑zY��I4Զ�� ���yt6�A�嘦�X�Ji��,}�u;	N��Y���@������G���n�h�{1C�uW�:�3 �n�"�����|%�jO=؝��ᮕ�lB۳kY�(�5t�q����r2���c��km��l��CDui6�nȌ�,���Nâ�X����fU�x�|~�b1q"��dj9K+�q�֚��]�����.�M�o��`�=X6O퀩��a���C����<C�DZ {J-'X�zУ�-a{���fm�7y���;�W��a��N#3�2��-�H� �:#b4��d��]�&���m$ �����7,�}RѮG�le;����:b�r[�����x[�۾�s�<'�m�zr!8��OOϾ�Ћ�$���,��u��l.�K@vر�)�(Ӭh�9�"��i�>$~t��G\�(��m<��i���L6��+��7�o�ޏ"�'R��%�Fʵ�2'����.��%y�c�f@f�+����]��I�Za�˿����|a��B�,��uCFƀ=OpJ�9�����cyT�RPP�Q���G��
Sٹ� �5���������n�0�o�����^*7���
B7
���)�/E�"���ȷ�ٶ�������
��kr�Y�^9�K�G{��_7�����N�]ԓ�]�׈���_�ݞ��Yn�R�;�N�`�����-������UE洛�#�ի�� �CeI���YY��ec~�{%j���~0\�!ٵ�P����Ŷ��YZ�ue�V΍��k��yOJ[�5����c�?~d��1��{l~~��N��U-倉�cƝA1rm�a�_�КY�I�#�\�mW�B���Ks9�ݘ_���Z�o�+:�+�dlA��A���'z��f���Ą���=��[���:�����ʹ�b�h7?&4�L���ܺ%����{(Ǳ\�L%�63��~���%�(0�7F@��i� �3 E���>�Z������c����"\����v��l ��l�Y2����$�'K��!W��$2a�s�6,�G���*��F�uE�q?���c8'��l�eO{��ޡ���i���@�ڎ�SW­/4m:�������(�ݜ�����?�,�m)�0�Fg7`t$�����8k���RE�>)d�<���d�hX��w�d�lh�̳�,�w��H�rr�����66�a]�;�����"�&�����P�x�rel"�H;�~`0'�8
��]�'}�l��b�\ݲ�"y�;�h�%�0K����k���A�e����^&�)@��F����غ�����*��#Ew.��D�n��|^r3����܆�%���A��H4�����$˾�{]뺺u͔�%�;�����y��?�Hմòi+���i۟�۹r"/!�o#���-W��c�����\�
�?��*��MmdOEpq|V:ۅ���j`��Wo �l��<���Xz���@k���-�6I�:�}
ģ$�[�`��"�?����á���c�S�c���T:�p?�H�(���j�xiG)��VJ^ۨj-���`��U���7�� .���)5X�~$��H���:�q�0'�s��Ɋ�M
2�%�{>&�*2gS�n�X����K��^Wo��д����=���t�O�����U�4Q�V��T|��W� kP���ԠUQ��������v�^^%AO	��K :Si�pr16�zk��^O��Ux���T-QO�*�-���	S�ɂ@#�>���R�ȟ�Ҹ���] �W�1JG��7ղ�X�甛�O�@�qW-8��}Ř���`Dޝ���ڜ��#\�1��r �ƣ�b�'Ѣ������kz�����������9���k�t��JjPn	<Q᯵!������l� YF�VOzn�[A�t�a։�J���ͣ��00��=Ór6�8��]�ٺ�{�U���Dƌ�B�����#��	K+m�;T¦����}.���WI�
@���(j,�!�>�x���]Q�쐮$�}�n�*:�-<�ȉj|4/A��0�UU�E�}c]�(F�u����9���T43����"��R�V8�KB�sߞi�伱�*d`Q��4cCDie ХBz̻C���$	]pf���Ow�Y��hd�[>読t�Ïf؟ڛ��l5O&����S!�<i���F������j�Ft�.Ύ%6'r\N�>	йpl�%I5�=]?Q�DC�'g�7>��C$$O���'����'�d'�����u���C�~����n�u���V�:��">b��.�\�vhB�vI�k<)���H���gqA9��m�M}U�l�i�����?�D׎�%Kڛ��rI�q�jYg+�n6��)��Q�O͂�}��0~����U����V�M�c~��"�����7�{�_�I(Z��U�^�sސ�\N�Y�_�Z�pkʧ�����piTF����]�U�sw0�*�A�F��I�`0%�*�r�|�K�ON6ˉB��WaT����Q��H�j�1�&�MK��OR�~a��Մ�W`^ц�I�mg�LN����
FV'�U0��{#����3`�Ϥ�s����Y�'؂��b`��������_�R�b����{�|]pJ�V���"f�X\�*ǁ���pp����ة�k��~-����l��w��#�
ǉ�:8��b���፷�9IҞ|�k>�#b��.�G�G�;@�jJ��J��Yf�F�|��m�r�"��ϐχkA����?ܡ���ƞ�p��� ������A�M����W�� W�
����ڊs�T���J����W[�S�>��]o�u��uA�O����\��ʏ�ѽ� �����uXr�d:�7����3����s�W
��������2x��
�˥�B�~`4�2+ѷ<���5ӓ|�Wu_a*�����i��Y;�>�e�+����H�R�f�`�pM�(�8_a�$M/�^E�[��-�(9s�ڻ�h�����k����9����.3jf'�E�h�ú �0F�z�J��i/g/����<]Rδm�ƺ{���
nO_�(_�*�qO�����{�� �?��0������B6��(�rvN�q�Ha���>l�ö��)ĥ�_�'��lڅf'�Sru�b~��r`���s���b�;�A�[�i��dlxƞ_漺,��.�~��ى89Ƃ���(�����xi*���،56��#9HJ�oUEc&M��-Tw���wŚ;H{j#Rk�Sos�ljz���҉��-��P���)ͨՈ�Ъ}ä���8d�@�J̝��BY�Z���,��E�π���(��+�zU�6���7݉oo�u����%�|�ׂ�^����4]7�mյKd�m�	 Ղp[�=G� ����{�p���}Dn��n��{�l����9ebގ��u5���]b�.>�|$���[i8���6�*Ihy�ݒC	���pS*�⩢,Y��*�����99��"����s'Ƃ��g.;Qo���ᶃUg��ߑ����n����������P��f�J�ڵr���2ê��=tCV���v��y�?�)��̵23?� �DG��}���_�`�u>}׻�df�=��0��� ?�AB�L��>�j�2I�]r�.��O�6���p��9})���0J���ڋ'�/���a��#M�J)��5��������6��-��>�:���2�>J9�N qU�O�*� �,�ݑ��Zܘx����b@��FA�n��x�0|��Ze��Ć�5�BNEl�-@��Y<�ӛۨjK��h_ˁ�JR|�[����������y<S��Q5E���Z�@��W��&^�*j-�;��$ѭ�]P�T8��� �,}e�D�
p-
�����E�����}�?*P��\�e���(��y�bM���gr�S܇-M����9��۫�t+=�$�!��cm���^*t��*'^����o�!�fD�V�	F̈���[�������oB[��Vr�$������ѭ���-awE��#zS�7$�J�I6W�dD6΅�5�5�/�&�(D&�5{g=�o�)T��@$��k��ˆ��� ȷ�;� L3(4�NYR�Ʒ*�8�;M�so@��x����1I���P�u�(/=?}����\E	����Ù�����Q�b0���v'�U�S7�ݚɇR+��z����e|I�^(椑
�/���S|b-�������� #�	#g0ǻ���N!L������4�H�`EkuH�����i����=���'G��a��H�S �j����R�^ύ=���]���v#�xۓ׊���M�%�b��g(�K����;���]u�M��9kIIfO*�B��?�6&�15�;�|k x<���/D*�B��V��;.�q��?Gl@Rbjf`U��ƭ�����ɪ;���b,���@��G�������5b�~��=�iz�+����ߌIU��N9�G����!����Y��ז�������$�O��g�����+�7��qcM'��Jb���j�nI�n�.oXn'��
�+��6�
����(Bj�	a��,�����'�@����LG����~����o��$M�U7pm��� �&0�țf��a��,_�}��G�cu��nc�I�	>��ۋ��{$Ymf#�p��h����jWx�U���_F�K�O���([��:��af�6d�s�7�|�+��Ђ���C�3��k>h{��Lᕿ�M�JD�sb:jv���6K+}V�}Ƚk�3.��>���8��>��px���*�$x�$&�#CW�)t�Y� ~D�����="4�!9�q��0�)_����������M�v��Q��2��5\�Gu&���y�F�-�s�~�Զ������ʫSfc�f��4��nO�UJ)��7�+��?18�)���X�n�| =�����W$�����l)K7�CR���/������[I$Z�H!��5�a6N��n�&s$1�$sPFL�l�H���ΝJq��b}����+)6ȪJx��_���l���#�
l̜Y���@�b�{	�����Xn5��_��S�O�����Z�s>�!�H��Z���A.�(�^V ������U}2j��hN;�[�3�'��Dk��e�RH֙�4"���Am/z�iJ��i��i:1!��&�$��X]LI�|B�GsK[�Y[�I��Uo��3O�YD��~_��~7�Va����0#%��\���4ȿ�38(�=�ۑ�(��k��Z�'c����U���t�HEۥA�!lb@�m0�M����A���	�\�Ѳ��by�{-�<_\�{ш��/,���Fi�V�X�R}��,���u�2��w��ƙCk6�1U�^[~;S�bK�/�d(�b�@�4�2��Y�P;�KC��Y=�����<�|��Q��Z8���Y��<
B.��K^��+�e��@�?����2�|�ۇt��E���t�X({����='���}"�Gm��55.a����YV���B*�/	.Ha��SdS�>��wdmmeK@�3�Ȩ��*x2R	����5qi҇�����9�����������z^ll��9�
��.�N�ׂY�O�a;8hZ˺2qZ��|Y(�y�݂������K0��0p��RW^�.L���s�N|���i���{��Ǩ]�-���M��,5��d�ѧ2��܇�1�\�lK�>W��Fۋ���3��i�8��q�܎ĚM��l����ȥ8ڄD��.I�]^$ .~�7m%�R�o��MbA��.D9Tl�z�����w�8ռ���A���!�2k9�)�ӫRd�j��גYU!|b�o-A�U����]�nR�<�{쀠
Uh���9������ᘉQ�]�V�����o�^@�/�~�	i9q�d�/�mR�?Ӱ�A�_6&:��ĬW�i��zC_�`��)i�k,���ϋS�Yp���k�x�#bc�E��t��å���S�W�K~���o�{F��X|[F�2�D��:^>w"{ݰ����j��gs�՜ɾNL96��5 pov2X\�D(��a��=��j�@���S}��0t�!�@/f�-�z�JI}�oh�_rk���',�,�P�ҹ!C�rW>�V9x>�pD.z�V�������Ϭ�ʳ=8Z���k���yx^�5��%���tj�d�u��9�i��T��	u~�٠
��,���Tf���@�}7J*�pȂe��A�4 ��#_�[���X(��] @��hG�_@a#�Tydeek��ǂ���� @8=_Hd0z�`�~��CK%/Y����3UZ�PNn!��ނ_���o<`L����e����P�(�u_�����D���2�*1m� �����>
�)�X���qO���l���h8�;��ˋ<��)
���'��b,�
 ���l��ݧ��~u2�6}kt^�
���t!uE�_)L�`��*JspR8{�iҘ��;�W�/6`�z���э��?Gɵ#��ɇ�o�����_+r�[K����*�g�r�^�i����+]��*m�U��Jg�~��%���g� R�b�
�r��o�jG��ͩ!Bj�hcu��}}�مq4pB��L�X!كG�����]@��7t�������\���|��kʖX	�hF ����N���I⡋
*����`)���E��o�������@L�è3Nf(�|�U��Dp��]���L����!���jY��.R��z���؛�9EK�J,���K�b`���Nqp�ElL��,�1��1����Gl��w6Z�x�i����$F�K�f{�:�v���9c���5^�p�;��|ay�d�������ԓ�&%e�B�]P�����nٸ��ԯU�܁s�o���o[0�`�b�����&3�g�agE2b�,�5ͅ5�]&�4��3��9,>��_9��W%��`dz��%'��|����o�
ꎍݝUx�ъ�8[X&��`�dG�v��9Z�����H7(/�w��c�CwX	�Hv1rv��G�T���qJȗl�rhr��\��櫈rz��NMJ��+9� 	��[�;ȩ�ll�_�6���:DX���B�޺@)�s�2���'>4�`�U��X9٩��l�u Õ�I��H���t��p*3�!RN��h�����O�V������4l5�7Q��W���T��Y�������Z$a����>-�4�G�w�z}ȍ��3$]���iE���C�E�� w�ga/,��Ě��V��#�j�z	�Pm�<����
:J�nd����$y/� *>�ﴓ�.��(�6��
s&o��^#�
�e3R�W�H@6��3J���b�����m�	�9@�c~�) z�ML���_w��+����F癮����r�Nb��;AH?z2��o�ۻ��l��N��@!��*�����9�I�Ϥ��.(�)��,}Bd����,�I�P^�;��DV9J������;�y�2^m�+���!:���$4���eId��GZ��G�kg����; ����_�-�.���F��KD�W���Ī���M� �15��B%:܍�Ǖ�r�4 [jٓw���A��d��K�A�����<��2BO�o��76�����K⻼7��Q�#³�l�=���:���Ȃ8�q�V����}�j[�kE��#��[ ߂��v�p`奒ց�����4k�s|�PP���GW&[��WG�ul����s�t��7�S|�3o�:��W�������ZؑՐ�=��S�6<�2�u�ӹQ���x��㳖��2w�B$�����q�!X��Ays�I0�x������<"�#��t�["��%z�	);��f4-$�$U��ψ,~|���0~B^ i\��I�X�!@�(��V����v{��P �ܣ<����
�M���z]��=�g�K�:��?�O��_���zz-�&D�=Ȗ��}j}|�U���;��n�MY��hL�f�k4����@@,�.V;��4�2�:�O\���k�D����.M�jF ً�C��]��!�67��Eu��d>ꢬ�N�A$j�!�E�|L�'��M��e�N���,��a��0��<���@B�8���D���ZJ�@)\/"zX3����k�Y�K�������"��n�����z���frSlӢ��)&��=ͪLg3)� ?���1�K�R�Ϯa���CZ����t�`���B�����ɵ��}���rҬH����efk��;��q�z��I3�6�˝˅k�n�]������ZU�0_�Ǝf<z�ޢ���ws�&6$�@(p��29�6��q��Z>�H@�V�)x��w)h0��2vZj3�K#��t�����2�p���?��׺-��l���逃uW�և��}�������)9��/��B�j/^��]�w1%ǟC���%сAP�4�̵��`ڞfG���m�D�	2!�J�A�t���(w$]?��)��F������V�~<4p�e�5�b�/g�=�u�;�����#>����4���٧����%_��ww����)���@� `Lb�Tn�&N^m����;N�ZT���p���ۖ���W���p�P�.���v�p�T&'���I�z�b�7=�t����?;�(�YO�5�j����4�D�0����+n����.���{��������A��7w#��+ȒO$��ߒ�4X�*�k�vi	p�Ӈ�PFz�L�R����YLT���=�9yB/�����̯&��;��m���:��c��W��	Ё\kٓ_�
c7��s���P���a���C"��F*�/hF��������ףB��L���S�JNc4�_�xq�{]y�͝��ٽ�L7�35��q��U�f��lo�ț��d�9AeN�����/��Bb�%���.�v^�X�ǻ(��B�ʠ������y��J@�����c:t�@�������Z>��1��J&�����r  �v ���y_�\hm���
�5�o��3h�R|��$?�e�67�d�X���y���ۈ�{U���@��<���̘N�|+���$��j8Vr���n����Ye���.�-߈L��4a�}I��;VK�y�y[.�N:R2E`�/�_�	_^f�K�9ty����3����o�RY8��*_A��,�W8��D3 ���K�NҺ˄�RyL�Fw��Gȇ*��������� s�[��F�$��0:lZb���^_�~v�?���8xƱ8�����9��y��^Kb��6u	�ǋ���@�eCa����4��G*٘Ҙ����1��v �z��7��g���n�v��j/��;`�IyUJ�n��ki���������+696�T>��dG��ﾮ{��&�?; 0=LϤ�=�.x_��Gy$�JQ�ʳ��D�%=W����V���7Ŀ��oƈ��KZ���ĶQB�!dJ)�p֏��P�����^��������h����j�������F<���}3�8#dx��K�7e99�d�G�la�+/�qs:�p}��A�U��>�"�0�34�y�Pb��T��>���펔P�a�os���34�&�E��p�bW�u?��Jy;Z�)�ᑏ�I�$;�d�����1ډ�A:L>ձ���ȀEc�4�����e��ͱs�׀w{�^%�^K���W;!ȹ�k�F�:��M�0���Z�,	��,/���'/���x*ʘ�lF�������1_�6��Ģ�W�q�ى���ȱ�̖w����O������U���l��+oarM�z�A��y��33�'���!�+3�q��Gɂ
V}�LӀ%�1�G%��kJ����Pւ�d�&�n�%����b��������0�d)�
!Ο��b�-�}�����S��H%X�O��,`��|�ٻ���1s�g:ޫ��1O��*_�]=dM�=�Ě\V*���˰M���;^)�6�ʅ�Z�#����V��e�ڡl���H���՟��Mr�OTwܥ%K� ���=#ks�V��F��!xk�Lc��Q=_pS����%T4Ǿv��yc�U�#Q�r����K�N���4�ޏ��f��a?��Fa��^�Xt�� TB�k\�bo�rʆ"o���b?�oDtLӎS���?��[�3ԱSdh����'�
��X�]��_$}a�d$��}L��`��c��$�b��񲀉�VkƤ�kDW���9B�.�|>���-sj�7��E�f2rv�+���:�E�\=T���jPh��!��� ������a|���K�n�܌��C�iH���'�7̈́Ft��N����gB���j���ȩNUbo�3��:�)#��Y�  ���~��<�n'4m���9ڹ.af�|;��@^|{f]5O)�|�U@yb�]���/��= �"��s��!��Y'Xˈ[jj�,���_�'s8lc��-	e�Bm�Z^�+���/|��wb{�:]�����nn��B0v�C�El3���J�(��|�Lǌ4B ����I7|n�gX���`? zzc-7G9�)߿0Ǟ����#2Rf���^���:��Э�
����*uM�S�!A�>䯌j�=�IF�D�:�[��U+Q"�-#Ya��[⫉qv@������^���y����9����`		�f:W�h��f˻�)A]*�>�A�ޑ�����.�p�,�D�f�2��"ɫ#�_�4i���6vw�D(��	�t/�t�qp+�<bk3��ï���e{�3Z���zJ�A� s(�tW+n*S��C��K��!ʥ����Tjs�u�'�hiS	���g���H��~�!	�|�������N�	K��q
,�����}r~^לKJ��z/�rDN�n_kp�L��k� M�������x��4w:� �����@�r�����"m�so�ux7+��?0^wƃ8p��!���|N:u��45G�b��!1Fis��,![�Õ|\zQ�
,����K^�8r>;W�凨F!��*jS���Z�])�O�	�c��ջ�����w�~*q���#��&�x��L�i84U+�у#�U�5q�5?)�d����|���𧇫�	��:�5����R�`�5gg�!(�׮;[}����PιY*���̲z���o��wJz'�h���Z=Զ"0Da�{!�~	�ҁ�cD-��I��ߊ��ҳ�����<F��Ǭ4���E�5�7�C��������/3�����v�i�P�>��f]gx�jP��x�-_	�2|���/,bSb<:޻� ̀��Y� ��4)azm
��B��C��D��:�Wdy�cB�����3�f�̪����ca����V�e�m�"G�^N�/��W��W��gj�ڍNPr:�v6m�)�ۨJ�I����8�0�ULbvxbߑa"e�p5=׼�؉�O����g��pi����G�Q�R���Su(����:V> 쯲{�w��P����+�:�Mz�M����<@�2Vz���z�9J�5D�Ķ�����f�N�!�Y?Q�3ǩ2t��X�n�ij͑���Vq���=��p����"Z+)�TěAp�O�����*#���6�6������#ؠ �ׇ�K������{�BR��l�>���d+�.ws#�w��������v�B��A��|g[O�C����*Pg�d���O+���W���fT�	��z��Ҿ��a�������=���p;~C�s��O���2���Ɯn�U�ުF����v.��4K%y|P����vy��>�k�u5�@-�6*,)��:������!;���c�c�sb9�������O��lb�o�L�K�y��7w�v������h�>��CiG]Zd��?�x|���z��Ӏg�ߙFp�V�	pԁ{e���	z`Ϊ��a��b_,�������HX�P�Oh�m�|48M�+��tU�C�!�VpJ2�0������:�c�=�db_gء�#A"��=f��R?�*�^�����vy/<��x��!��.%�$"�;����"�ꬫ>�C����C�����Z�zc�js��t��b�^l+�m�i�~>~K����
�;��;��z:�kO��f�v����F,�R�蔋e�hU��pe�6V�������M�@[��Ϟ.?<|��-5���o�	+<�ݔn�&��H>]�x��7�׏�Z�>�F�G5<�\��\/�"<�C�����%��q��q�:SL��	|�3}�܏�<B#-8��5�j��`[�p��[@���N��1�#R�a$��F�&.aNv^O)i]�>m4�x�����A;C1I-*#,y�Z��8g]�P�Р4��ү�(@���Ԅ�7�h\_�Z��iX����]À����6�������<Բh	�����^0py�Սp�]�Q>��?�5�"��0}a�>uwY>����p`�
�=��+qth���H�, �7�m�՜�9L��:���IJ=���5�ip�>ɹr�ڠ|I��tW��8�1��Z�XH{�6��eǁ��詇3���/��F��������	��w|�G�4}n���?���l�g@]��
T�SMҎ9(�U�c̀@��Za~_�24�%H��l7�u�?e9c�d�FT���n'?���_�U�i�r�B'�<�%.O �Ŷoi�k9_�g���G�r�i��"8�)_7�gTO�f+L?��p��;�5�4��W����'�8��N��S>Q�=����'�{W���>|��If�[X�8>F�K~��R�ޞ���Q��S�+�"�����@��� ��Y���
[��zq)ؽ�l��&�u �ltP���Ԥқa��J�(�G����΢ih��	O�Q����a��z�CI����`��ܢP�w����Ѣ���JmB����=8�>�l&�~�Dn|��V����s�I.h�ď���A
�a�6��,9����"z�������g��11�)�e��OO8��H��w�Tr]P��|C��IZ�����B<�� M��I+���C�}���3����j���B{�����v�>�a����aY�p#��b�'	!R�
�6�#88ד�P!�L36Y�/�5���ts���Br����.���&��#o
3*t��RO�F��]����b2!������J�����N]�?+�H���8n�1��Ual�ƌ��N�+�s�^+^Z��������[��&IN���z=}���Ǫ�ߵ������O�߻��p�A瀴k�&a���� s�"���%EJ7�;�{��T	��>�CfM�4X:�@�b��w��{�K�4��J[O��.9�H�^�5������S��]�;5���:�4�N[5-,��OL��s��u�Gf���lY;�5B�����`j�fxaVv�`2wӌ�O��P��橷$ �1��F�5l��f�iw�A^����6�	�H�St�X�|�HO6|���k��DJ=v�ه��� Zaċw���v�s�����%*�QnQIN+nI���G����!��+n"LW�il"V��EI�I致z�`�V�̦����0PY�7�R߷Hݨ���
-��L���g&P���Rz�lsj�	`ch�
�7Q#�)��,��T�Y��7�@���5M�+_\�ɛ4�K��ޏ����ѧ���:d�P��{�pC"�p�8/,��H�p��/kiYԒ<3T�a�D���2��8e���Y��G���Y�lѧ�/7>��ȫ1��&XM�D���i�w�N4:��P�U{5쾣�����V��f���'�m跁��|5C5�<eb�Ox�뿝G���m��<\�)�DIt�0&����.a<I���bcls2�A2%�9^��*�"�#�_'�'ʖ�A���bPq>B�@o�Æ]���X�brw��?[W�%�FŽ9 ��v2؉)� y����b��9��k�0P�R}�^,��[Z/�$�vo6� �uf�'�c���x)�Q֭�I(��P2�����r��j��,�0̨�s+���lW!��Ml������[li��t���5_��X�ȻA�/x3sM�-�F����%/�i����J���aj��ʋc�����MTא�͔�)�T#�K��߽Z[�r�q]��ϰ��g���%T(XW1IV$=�g�b��~�#�`ɲ����T���`�n�B>;@d�"]n�݂�C�K�FS��b�kX(;n����G� ��
P�3$OOv�(��c�
�y?$ �S[L�I�9!��4�`�t���9��L;/q��3~Ӭ��LS�C��m�]�n庲:���č Lu%�|��6'�yW���s���p�q��CZ��[�>Qy�p-���
;ӳ?�+3n3Ν�X\g�I��5e��X܊#h�\B�e�gФ��橡WW��>��(�*H�<0��AhC��g���|3%i�
��v�6�k�zE>؀_��b4����[&[_4���eOh��� ՅA�#D��fvI�cV$�2l���g�������a��\]X F�C�,I��@_���_A�O��ŸB-n���Vr��Oa�۫���Q�c:kA���-�_p����̍71�!���� �$*V�%Aɥ9	+�,���r�x	M��mv%a �x���̍��T��%�1�6�Ps�|zB��zw��_Ү���?C|�&5ڙ�BK�a�Z]�������r��B_2@Y��L��"�Ē�yP]R�4d�PM��U���Ũ�Jp�mO�c�*@c[� �4�p���0� ��||+CG�)ܫ(t{��]��sGguC�|��[�F+WƜ96u���%k����6+����F�S���k���y<�$Tf����76�)7�������Ŕ���B�X�"`FQ��(�	���$�=5�ř��0S_Z�4 �a�N2����ٴF��2�+s��^/OWKe��9�"ˬ�rצ~R��e��YJzv�<D���U:ج)�!��a!S�f�λM4�ۙ��2NE���E��i��RP1_�c�2b�i�Xڲ�P��~e�ԠQO_���뽍�ՠ�m��6Oﻩ%ʝA(���w������A�ۯ��`]�-4P�m���%d8M��/Ѹ�
BD��c}�3V��j��pF��^v�P�c�U����@& '�0\�a����f��GB>τ��M�W͌c�ƽ�^ �'鉞s)

�*0᫱yJ�c�a������Ň�v��o%�\�~5�y{��y����ҵS��n$�<O�������bȉtґ*hv��e�g_+�s�}�� �e��9�������Y>-�7�KC�G��-J.߲��0,Jfڜ�m��yp�Bv#U��ҏ)����nh{��E���D#�ȭ�D~�j<'�����Lr�6�6LT�g��CW�Kr�yu��$�x���Y�����)�KC���yF�&TE���Ģl�Sq���-��PϮ�B��!�]�N��Ewt�v~�Ӱk8&1n��m�2%
����q�����[�cl����l��&n�	���J�z@���㌟�ՊfA��|�^�Xr���C�������|#�p��ϭ1Db�1Y:�7�l��:9�8�03�T���ތ���Z��9��1����
\�ݏ�������N^q��ῲ����D?�/.�2��0bT���>?Bs������Ƃ'B�r�k�3�;��� ��N�=��]t�sU�
��h����q�6��⩑f��홏%���ĵR�R��H(4g�(��˸���=b蠉O�͏���X
���C`C�B)�*V���!��8bxgDV#��eNj�@��}��/��Y�c����刁X�����D����xp�"a�&��:/o��`Ru+7�5f�q�&8�TB�.���cG^���T��=���~wí7�5q`��t��_y�j�Ⱥܿ;*;����؇7�����x���������N���7�>Z���q'��Ǐb��x{�i]�'�e�}z}D<ɽ���X��Vd��+�m�c�l;�N�/nz�p=ҹ#�S&+�C��n�(�l��"�y�z�DVs8(�����Mf�̽�ͿσmS��g�zQb� ��Q��\�φ ���?�L�}+�d�1���\�_N�[����	�]-v�-��݀�9�c��	�������/	L�;�PdHכ��(��.V\����.���5^��I!I@��e߆�M�za{������{9J�k�~̆�%+��5Rtv&�7K�P�*n��<_������e�NY�/�><����Ze����p��!�<��8w�1�:��נU�r6��Т�_�/� ��~#Ԭ.�T�	Պ�cp#B`r_��fC]������G���d������\M=���Q�&3��02@j@��-h����6����>���j��7{�,$�b{�2����m��~1d�����ZN�I���KzD#K���B�(�yn�K\��Wܛ��N}��W�n4�cdqQ��m�N�E�i��kҟ��Os]�+����{`��ˮ�*��q�<���f_Bo՚v稟��6e�X�V�cO�9���I�mܰ S�6��!�?�"P��"����u^Hx����D#��V*�	�2��o�jv�Eq��]0�U�sSUF�x�qw�N�AxJә�/��g�$��
�׽�P�_V @"�yx%�P]�����&��ޭa:s�[M�v���"pF� YR]s��)�����4Y0��`�FQ���Ԭ-/L��EΚ�ü;����̑y��㑣���#��5����E�],d��F��C��v1��=ש��A�#A�.۰�@c#��I�
�w���� ���%����8�x�]�5�V��.�~����y�t��,�FU;!�?䆲(�+�o}���\�7x���eU)�?�S�������N��dh�cN���b�֐s_��O��&�)��m"�ʮ䟛�T9�$��蜞E���;��׷��lc�́��i��1�N�7����ª	V��rV�����v?&+.B��J���$39A5@����i8�bf9�©Q�S�o���!S��`pߧeOc-\>{��虌Q�&�.'�{�+q"�;.O���Y_*�h���#]��\/L��M���⪤����Ԏ���L��w;��E��A;��g����]/\ݥ��b���vIS
u����\M	ӹ�eǡ�q�j��K&�0�!x�`h��5��N��iJY�7��E�3`O�*�|�Y�D���/(�D�u���g���I�F��������\���3����B�'�������c4�zI/��Բ�I���cw�����$��0���}�����Ԗ�z�J�H���k�ɭ{6�BF�����>�S�Ȁ���޹7��h�L��%��6}@b��*�;�C�݉RwW~�J$�y���I���n��K�qD:1�s��u9��WE��\(Jc�y2R�φ��?��IN.��V#"I讇O;P�&ᱷ�_:�6%���©J��!R�1��v�E���ȫ�ѳ��L�,����Ul���Oӷ��@
�ߦ:oa"�-e$�7-�JMu{Z���`Q�*�/fL�c�G���"�f�#����6*��)@�h�C��@��6��k�/�	O�SP��q��[n�X�u �����g��$�b��u�(v�� ���ĕԭ&�s�Ơ�bB��v�kYʔZ�O8,O��`�?�޾k!�f�s�M̓W �y�)��`��A�7A��=6�����I@����(�~�Q[������}��V��zm,d�a�sX����5lI��7P�՟s��kY��q��_�!EP%
�o{�̄����DgQ������v��I�U8%i%5x�U��A.B D��t��J����1��+��ĳ1��yA��mK�:r��	���R���?ܷ�XL�TQ���sX�Y���X��;��E.���LWٶ�b�v��z�IF�sT�<�ey���R�V=��fon�C}~���� O��؁H�eBZ��|
>sz���$�&e�$�p~� ��~������@���P>�&���ϡ����~��k�ԍ@�(;\fXY�1lGK�[�!�,���ƅ�4w�_E��[����TŚe��p?��;�=j�����+��(4ľ;�qBA�f)�`�F!�3�a ���c�I�O>���:_`B$��������n��Tt���>��_�{��Fܱp&F�w�6�=��d�_+?��5�h[�[|K�s�2 ��"�/}� ���v�Q��wS�'�.a�Q�k;^W
Ǯ�6�>�)m��ʱ֪��9͞������޾;�5�����g��0���q|ꄟ����o?��9e�,��;h��jN�YpŊ�0­�W�1vs~@� �䑢g��6�tp_�2��c�I� H��e41)V�Í���ִ2"cf7]O�K�~`X��Z�Lq���O�;�zE.:qM��lH��EmE1��8��q{�� 㛝\���� C��y���v�%�,1�&
IŸ��+��|Px[:��p�Mw�T�:��c`_�Z���� �k�꜊A�( 6��r\�̬1�[\�́b������d�獗1`Wʙ��}_6����)�*�Q��̱z�ǁ�	`�MR��^�%���J�*U��)��e���[�po���U&W�P ���^$�37D�����@X��OH�?N)d�q����zbB��@���PM�Mh�`b��,�8�;���) �8s���m�]@� �EP�8�ҐM0.D��^�����_ت ;k�{�W�a[�����h�I�&ӟn�z�{�5�G�&�c�Yi������U� ������oC�����r�?�r|@A�jO��"\c�z,eFx���U��ua	cg�
������Y���I�e���͜�r�l>`/Hc=D�d� RR��o ����,�: ެ���̢g���&-�P,�-�#� ����w�/3��λ|���w���T՟���R�����C
ZoBF��*�H���fө��f���0�"��)�!�@�$�����ꊪd�2�t�7���Oڅ0���wѾ[�Yz�3О �K�.��2%�g��tqT�ʶ�5�q��5�1�p�炴��o�u���O-�_���'x��Nw���K?�8q�h�ĞM0{׷,�	�;&�S�X��W�z3 ��؃�M�����CzݦlA5���&ä9?b��";i���X���x{���<�� ?I����4C$�_冲m8���T��G`��z�_� ��@x����ڸ:r�'n�Z�X>Z��>��V��Wf��L>�J/��2�y"�ܘ�T�VCsQTQ+\�}bB�S��3_`Cv��-��NПqR�ݺ����V�U#�tg��~~*J>=UּaO2�D�U�Q�&���=z���P5�5i)�x�Յ�Br��T߿%2N�^���K
�ȿ�h���4B2Qvqd�v~r�`���m��1�>aK�������ʗ��p!�Ǧ7�8����]�oA?�wLA	��5J�>o�a�2Td�AP4��������O�]��d����jEF�;�Ц� G��U+]�9��]06�}�9�W�G���Knk7�l��AnPebX������}�ƕ�8Hq¨E!s<�'�<{w��x\������l�\�����_���>�ϯ8R�W ���۸pm ~/���e�ku)�OD��oQpKa2��"�ܜU�����ڌ�����X������n������n��$���F��/�e�ʊ${�~.Ԫl��~����o��P�QI+�6�̖�w;Nf�Q�F�_q=���Ϊ^1���겜��ga��'�3G������?�PC��:w�=>�(��P��4���	v̛�A�u�=���9VX-�u��6n�C���8�D����<>� s�V���!�4(W��Ӭ �w�����B_/�:�$Z��^>g\�8��Zp7iG�4���U�R����n��ri������С�����c�E�/����R�-�y���T<	�mGa�������2J���֦��d�$��(��	���6��>1����ccj�j���n]����5�����;���BQ��e�N�)�Y4�w2!E2k��
���n<�	��k��5]��wd�|r���m�����:~"a3�K��+6DM��;j	Pg,�8A��/�Eȉ�p2����.|~m�YΛ�/퓬��KJ��K�6B����	�U��H���VI�	!�*��o\��<�Z2��5�{r<��x1�[��}��������T��՚v��K�k�"�=6ղ�0+�*),��~��7�tk�s>i�H��m�11(;��S�-�VaY�`zcʋ�Z��`�ά��I<���J��f��~*(�~[�D���,&�K��X�1N��-_�H>.���S-}=�����4]Ʋ���ԅz)���E	9��<��u�2�l�ǁ�m0u�-�Q�r�������s�0�}�(!#e�ː�k�@��SC5�z �h��1YƆ٬��V����?�]w��y���(YKT6���1�\����miR��D�!1�]{�7���Q���ϊ'�3��۱���ߘ�=o'�����n&�Np�PB�?^���1�>�ϘgO��v�|h� =��g������������ݺ���x�.��3?5H��6���Zu8�����b��5�U?f��-,����;*��qa��L9�ϸ�aP$38\}:N`#=no3s����}�R�ATD���֔>ǃ	�����S�no�@��W`�@ҎȊ"�Q�4ê��1�uH�80�P�q���Դ&���b�O�i�R8.�e�b~ϳ���d+L
MY}a��s���B�[�?�b�9�`H�,�L�%OURC~6p^;��R�:/��Mk���n/Y!��OO]����a^T+�$�:,&ELSY�4v:�Ou%Y���6���mu�U���CX��Y�G�'���o� j8f���Hy�M��Ѓ������e���9�_��{gV�Q�,yB� ����<��p%`���2(��,q�yv>0�#�v�`7����rN~�BX�}�N5"1�����z���<�nd��Wj#��гʲ]c�9�F���(�y͆�0�yɿ�a�=��Fق�ѓxA���{����{唺R�S��Q�5J��,�$�����J�b�D/�sk�����Tz˭%?�`z���`Y�ѻ��29gJ6IN��R=Ϸ��1�>���aeUހ�B�\�Կ���V��R���Q����Z��+���7��P)Fh���C�9d�WPd�s�	�N��-�,�Z��.��[���$��p'F��#OO.���06+��B�*�$D�$1�k+}�`P��FT��0��8��e�Zs���mq�&O<��/i�z�bQQz����RFfD��6���w�[p���M��bX��^�l=%=9q�k���KI����;�()�0A)�e� �AG�@���SQx���XYgm��4xK�p��v^�����n�b>�i�i�����|j�޵����=�> ��|]�J�w�=z�Q �3Ho.�D������p~��g>n�>.�1��}5��8\��x̯�6���M'ƙ�p$�߫-X�շ}�5���a�֢b��w���\W�9��K�}��NT�7b�D���$��Nۄ�Q�|��ふ?�bUY�?�����(�cFH�3������|�%4Q:���"��:X�~��3� j�T7wunGû�&�4{�jt�(u�6{�y��l�Ϟ�"�ظ�u#�S&���0>������jo�����0JQ<���)����,��b��o�����6U�~e�����`��?�7=��qZI�eq��������p�U�����YT$�xZc��S_�a�!ުٟ�Δ���	�M2u�f6�MI�I��2^��0�Z����I?^���2>���P,�TK�ʩ�%����^���w_�Ix��f�a*�X�*i����\?cf��T�xQ0AH8�q$��g�$�p4��d2D΍��x=پ	q����r�<]N�����n,V�����pi}�3�#.����-,�'���ҝ�5ˏ-"��� לܹ���*~^Z�/7ZJ�0*�V�>�E�O�@q�	��6N���c��Zhǿ4�!Ӻ$4��cm��h]>�Ƒ�By�NA-����.����`bV���t ù�-/ȺX�PӠ�s����d:�D�H��$�)�U,����dPF����u|;?<�j�+�Ec@4M�`+�@��A^���-'�������
�q�Gc����c��`%bUOgH�W�?��<�ȿ8�rZ"���̞�^h�L��>B9���R�`��Q��cxI�9�.I������wn�}�[C߁�;���k�v^�i����Մ��D�X�N1���?p�wN�s	0`�z���Cr"��<�y� �x��H�WG�_ �w�����!�}MҎ�� Ι#W�&`pC�А����Ӟ_�<lM%,x��cƲ+\V��r�{� ��@�o$f.;���C8|J*G^����?L��$���Ŕ�D���� ����-��NdgW}� �eD��l���?�O�q�����.	�g	�h�3^��.])À���-������ �E!h�HW��G]hխ�E������8,G�!s�e,��۩b�מ4�����1<tv5r8=�UJ�\m�ȅh[�xvP�y��	Ur�c+Q(�T,k�vl{�pl�"��r�k�P�(�S�!�V�iߴ�W�{UM�d��d�dM�0k��E*R���Q�b�C@�X��1� �B���cD@G�H'��zQ��_V�˺�V�DD��4�R�ԧ����k��,rϗֽ�qj��l;����=N)*�)�w��V�8�\�ޒA`��G���[�",z��
�/	�g�-_bɀ�d�s.��FiYN$�U.e��n�.ĔT���
L�G.��S�$�/�����D��$��u� OkB�f^%?��)#|�Ѝ�*�/��K0}mT�[�X;BK�[�ը(��4Q��m.�x�ܔ9S���ܡH�D6a$�4Յ�N�c���:N�!M ��m�_�=�)�)�蒊[�`Tݘ��QZB���V�;[8�?y�����A�͊Z-��:s�����e�g�^�:!%3�?X��%c�/��mN�ip���:*���lB����K���9���L�6u����\�N�?��,s4O��I'�Wp��p;��;�EJ�f�{���K�ej���<��;�DQ���+>�����!i���R�ꅶ��K��L�ǆ��`����@�aw���d L�6p��|��߾ȻH��`� �2���4,i���V�v)t���Y9��F��C�;RT�w=.?����g�+G`S�����Ma����O�̧�q��P���ed�	��H�=,d)���J��|4b0��6��v\_�n��Z���]�h�^�2(��PI%y@�lZ #T�P��c�mvM��j�T�c<�t���������!6�����u�)����M7uvt�ת�Pɿ/G���Ԧ����B
kB;�3��`�uGcl�A�H4$2�Ś�N2���(����0BI�.F�H62KQ0,'���&Ap��?pSdZ: ���z��ǹd��*q�s,�gl�2�n֧~�,6ۖ�4fQZ ���P<;z3k�M�4<�w�&!c�q��J��q �Y(ȹ�:-��{��z楷�ŀ��S�&�g�qϚ�T&��$���B꘎7�������m�	(��⬫jP��{�4a	���Ɨ�ߖ<>�9n��H�a�X/	Q���as�-��Əw��/p��T�A(8wRͅ�ݏ�EB�t 6�%�j�A�U�Igr�(�/��q��-cw��F��ed(��?6R�A-���e[�� ˇ� l5]�񯩺笨?v��ݟ�.��X� �%%L�!�����
KT�.u�A�ݣ��*�|NEt'B������He7M�	���� ��|��?D8�o��(aQ�}R+�Z3+�V}Ǳ'sf�ar���ӷ�
6	���&w�K����>]�S� �����e;ⰧE��ă:��ݽ�,�R3"s'pR��H����VD`J;����۶��v���6��O��EUYP��f��|�Z�m�4�q���3�n���Ã�h���.Wf�{Jf�ۗ�:��߁f��}@��~_�t휩	�`��bѝ�v���������w��r����R�������-?:t���gT@-�0�����\�,^�O�ET�'R��U�ax�
�`s�G���u5� ��7Δ��LSkޛ]9;��9%|��.�`K�uK�Ω�tx Ϟxۥ�<�Đ-��8R�
`��4�Y���ƾ�����5��BO���`�YG�@���r�Y%���;���n��d��:�NR?[��桎��'�Dņ��17d4'�����u$�)�c���	l��
%����7��:l��q�|�<�U�P F?H�r�����)��ϠԞ[�Zٞ�����+D/�;�0|Z�`��Hf���~コk��4Tzz2JRl�A��g�n?��$���+�xCgy����bV�U�L��{v��gYS���uҽ�b�8��H�V��-
ֈ����S
j��|n���Kq��p�.#��?��Μ���R�$������b�SٷJq\�bh����k��E�ߩOV�)�1n�<���C�̟$��[�����ek��#M:2�U1`:����x�׏��&~�;��+O��;�;���eL��|Vdh,�����%]7T"���`�^��J�ʃ���k�ߧ�_1�岹,�,10'�sS����z�Ip��k�b�j&[�Z��F�K+h�#���!c�>�ɂ����%zJ�|��]��^དྷ��q�CѰ�t"[(:%�b�y�5��gs���h�#^z���P`�m�.\z��)?Fj��9��)&,��q�j���x㽖�;Z��ͳt�����O������~�,�x��6�>\_�o�<vҋ���2u$O��ف���{4/'U����F!�\�Ys�ssy��#���Nк�,�۽Y<"r�"Cx���,\��Q��\�x7�PE��G��Si�υ���H�D�X(���|a�%6}�����qdQz��/3��3����Bc9��AAE]��	�s>?�]���Z����Q��^�y���5���x2mF��;����\�R���~�7��ai�_,s��Ǒ��֡�ꯂ�XZ��U]���~�hף���9�k��|f� @oS�-�U���{c��������������ͯ���s��;¨O��͕}\�n@�P�!�N��[���F���*�hk��˜���$7��Җ�,:r�6�3<sE�)t}�F7�Z����^���L�.��0�z�fJ,������d��qA�^o��c 
���+�������u�@���Z ��--�a%���޹'��)��\�p�r�s��A��v{���C(2l1���P����Z���j�^��K���g�G��?)�/,1L�|n����iÆ;��M���P,�eU�O�F^�v�7���J�V�U�[�=	�]	=���o��J��]EC�~T�A4����,^��z��k�D���	L�@!K��u16�e��;�pgWd�w�8Z�>����dQ�`m��d�)�D�w(@({�$)�<G��v�9F��!��~Aq�u!��_ |��⒩�)湂Q&�?���lZ�s��/�J�E9��>��ӂ �:�:��cP^N��F�jbn���@s���]���go-�c-��aDJ�D3�q�9,܇4P��"�����-H�B�ҭ��?��,�T��>��
P}��;���:b��M�.{��a�����g����7���xa�\#�,����mN��?�4]�	 �J�W����qn�!�50�U�:����F����+6E�hK��gPBC<<ĸ2V(��Y&ϭils���7����Ŵ�'�cB(댡t)v|�nSZ��R�ųpn��2�eȌ/@,�u��*7��H���BU�5)��%)«w�_��H��s���|s��U���i?�^Y\��w�n��SQ�U������fj���>a��O���	�𤑇y�%������$�c9������V!x��`I�8��������%'/-^{
���h�p{�MMݮ��ީ;k�w�K���������ф��;_k|%�����1�圌:��0���"(��k�|�����i�n������9���h}��<��T�1Xߧ$�~���@<�a��f}:g��>=DBJ�^L֨�ź�L5M���	�k�a�=6�ΡA�MZ�.,M]�@� �G٠�K�����.u.��&l�	&��n�����u�I_
-P"X���#�jh�����s-�tz&g�v����s^���.TEtǣ��MOH�2/=5ǥ�ٞ*���S� F8���l8m�a�z�ƛ�Uu9_լy��!aw)�ghϳؠ���V+b�^ԑ�����D�o;��"Q��{�%,%a����
�����0I���l�$��cQ��a0�y��e.5�q��,5m�84�)�ڇ=��J�5@��p�D��\���59�Jw�r	+����O�{��W�@oAnש�R���[Km�_�������:O��u:ᅍ.���Sw#��]eăϧ<G�-�Qo3!J$f����N����n�,��{�s")\�zr B�������G}��������ȥ~%_�f���9����ȏ#naCJ��ɨs֧f֖o��9s{kPS4BȘAj%p�kq�A�]���$4�a�:~� @7n�,U���{�G7��CAxo�hn�d���X��'�TA3:;VZryui*׃����)J�'��8
b�]�c\��ˀ�I<�{m�����k�f��j\��-I?c�rB\���?�0O�7��Eڳ��n;-p�	�Xl�3��aH)cz�G�
�o|�Q�8���NѱH>ɂ����zu�ݽF����� I-DP�-��U�|}��7��j�,�̧
/�����;֫p��2Đ/B�?�O���B�u��Īz\������%�z2%"�=�5���*.ch���������?È}2���;ɲ;�6y��
��CI�����{F7�y	{G"]�'@fbR�$\r	�A:H��Wy�o�r�~���_JL��1��]tɘ�1(#���������!'��4���ǋ�|�`3�=2g�&n�0*�=�:��Xe���N�΁�c���<�y�3P��t�y���<m�ӵՐ�˳�� Z��d"�p�)���bp�2�:Z����A�d��q���r���e[�����j��+4��5X=F��_��7W
D�9��g���&�����c��F$�m�s�F0%��M�������~�A�ii�%F��i%G6����s�{13�(������3�� ,H%��[#F%�ʳ2�]I�>$Hv �%]Ya��y��4�g���(,@e{�^�?h�'��ӵ*�${b\�֊y2d#�����
x��	smh	8b�D���W�aˤ�S~$*~��K��5*A���Z*�6�K�Ng@'/�a���_��I����,��dZ|	Ƨ.���!��`��.&����

������1%[�s�-R(�-^*������%$R_���"��s�@4"������������F�B���&��Fc�Iq%k�k��C����Aīf�[�Y����f2�V�Qf�U�ZST��ոKZ$K���<볰�mz-1"{��+���������m��D6/��ϝ
W%��L��!Q�*����h9����X:}���+��&�o�`���2���G����b#, �ן7�׈�D����!#�֧��J،��Q�G��b�T���}c�rŌ�.yD��������O]�#bqԳ�RI/@���"{x���٪� 
�����t�uH�_�a�}������9��; w|�Z!>����+��^�Ԅ���:�3������ݺR����.!xl����&�IqD3.����M���N?�`N�f���Z�}��_qZ�8CAU�.K�K���6�Mu�vw��b�'};py�	<���_�xĚ�@L��b�"�p����}��c��y��ص��z=j���b}g?��vg�A�:;O/�[�B�>���G�S����R�rڈ��R�>��C'�4�vbîS֗7��+�}I���dR�r�"��蒰��KE��q���c��jO�+S��� �:(}�#Ȩ6��2 ��,�jS7R���y�PX'�%���휿﷮j|蠲s�J��o�B�Æ�g��	����G�]����#��~�=� Kg���N�W�S�n�ڈ[��j�LE�1/��W�H�� �7��A��k����q��|O���N;�vO�^Yc�^� �ʦ��'ˑ<�́UD�ڪ٣M�j���G�N_�	���1�/,�L�Q�����T/�^����
�$Q����Z�%��qE�
uwTp�x�W:�/$���U��XQ�ׇ	�P�9)!y#4��dbhuUᦋl��.�M�%��J­���.ٔw���s��k�c)�� �+o���O����R�jNʄ�[ו>�j�!�����ڣK�*c�\ߒ1�\.��G���jxzu�~b�)�3��|Rj����� �Ab�K��R�Y���&v� ����	n���cs��d��y��_�)9�̇��K�֋�}_�� �D�I	NYZ��r�LEI�åg,��#m�La�h�p(?U ���d,n��mn�]�ƈ����/�[%����D�
u�,UO]Q��\+	�y>n:�c�Ǝ�զPo\�Yv�l�w�`����5ԛ���/���~���n~c4���5N�F��ܯ�>"l><�>w�"0=W��h��D�H��� �hW�&�q2YTIT�j�1�')W<1&^�Z��x6��F�J���0!-�eV�鶙�ހlf�gM��7��:9i 	e��ȕک�� �f��s��*n�yQH�;V�k L���E<g��t�.M������1�\��	�0M"��b�:�.��p�� �a�ٳ�!JqAb�M+e�prd��UO �X�A���fL�n�� �ۺ����5������60���\Du����(z-1*W��}mı�j�c|u��0��P`�ǝ�7��q��u�@�������'̄�����bdY���߫=����&�~�~)v*����óٻ'�O�8�<`rN+�z�_�K�"�?���	����Xuϑ�B�R���� �2?�P�/ӿ�g��}��S{��j�����G�
�v���Â	c8W�I���<v�`y�Ԕ����M��5��e^9��O��t�9����@�&�0�R��'-���h3��:J��n�ctF;s��w@7'�"�{5��	��3kG�~^��R�5b��3Xi�\ @��:�1?y�[�r���s���f6�5~��F�?�(�Y���V�Q�֞�;�?��ߞIg;i���d&)6�l?�:�as%LKXῤ���]�t5�UR�����.��*�=�=n$��]�%|�����w<��L����i�)�sh���h�R�U��
p��������b��Z��Մ%�ct���4<t��uͷ��Uݖ�"���*�
�~v[�3.l�^-�T���P6=,��#�/���grhM}$3ι�Jb����f33�_z�w��%X)��T�b��x	����4o]K��Y�hңېUA2�-;G������4L�DcTG�I��1g�}--��\CP����p{1��#1wK9�����zh��<��CE����i�A��z������3��	T	�Ā�!�&������<�J�T����AO����C6���NZkuPp�7��5V�B2�T����H��& yo���(�qM=]U���7�2��{�w,S��Iw��\܆Nv��y��G�#`Z����>���t�˕5oޫh���/�	�n55e�S��ɟf�k�i��.�$�]�1/}��@��Q�e�a;�hkhD���ռ-���SR8�`=H5��T0�5]�詛/��O���9O[ŇCo���AZ�ε\mJ�9���l��c&��6C��#�>�6�{���>TD������D�HA��9���ˣ�2��K�u5c���aSƱ��s�{[���w��Ř�~� &υ�Ӑg�}�n����ɺ? ]A�K�p:�h9��?;�AΡ����8��i^��o�N��6F��zi�Q��z�"8�o�7�mT>��_��o����"��%1L�ჳ��-�j��4����Dj�^ |�h(V����2�6ߙY�^D�Z ���R[7�n���S���7��H΂-��u�&��[&
C���D�����s�·����rN���K��PϿ���"`+a�S�8�� @�ߕ�Ta}���Nr��6^c懛;e�"g�;���=�f٬E4T�o��L8�V.�_q _�KZ|���B� �f͉s��%ŝ@�;t�6��Z`ОA��Gf�J��F���[s�+�PݐZ��AV�j*�������}����#�>�����ACÐ�a�Ox�"B�C5�SPyx@�d������O�k��V��
��m&����.�/���Q�8����r,�	r��/��x!G�{�й���!��|-!N�cX(Տ*R
D�)X�),:,�XV�@ʎ����٤{������ЅL|}5���-4Ĺ�І[Wm����\=�}Z�޵`y��a.["v��h�O/��0�~�0�6G�\�ք$�g���z��oȦU����{��ƻ���"���Ϩ-e'�FP��w-�������R�qB�дTѴ=��=.?0��B-J��A4��E׿(������I�u��(���5��#��t�=nC�IZ���m�Vt�-k�$w�M��b�(���yp�c��-�G�iNSU��{9#N=Iŗ1���By�(�.�e�7�?�U���j��W(��N�6Kh4t<�A����q��hN���b2���7O�������+Es4���瓹^IЇc�l���-�e?�^��O7���A���=����!�h>lK��M��g9x������E!
��0�T�N�JA~;$-��<�P[���O��=u�^����
���}Ӑ[���Y7#W����RL���a��k�]_$�=ݨ_Q4�=cTO�DK"�/�]���hP�2�Y�a�Ry�*���Oz�pV��
�qE�}SuW
'o����#t�,����b�鞎0��/��c��:mF�ːe�py6��)��2���*f�n��#�o{%?�1I�
�ZK�qX��?p��%�nd�l�M9:��CMk�W��Qp*����L��)�ʥ�q���ғ�Rq�E�P��8�D�� Js��Y���M�������?�^�~���/�m�[�H1��j('	����ɨi�(߾���1s���Hhg���Q]brWiW:��N}�����/��PH˖T�sܷ�(�\[�/�\p��2����`ӿ�_���F�TK��+����!-5|��#�v�(�`P
D�����,��Icn���%���IC�&�:a�f�3�(q��|���XJ>�e�(��y:���a�n��O'I�.C�w���{-���;�H����ỳ�v�_k�<���t�pC��2O/֦Lm;ou�f@�g��V@"���f06��7y�N���2l�OxU��<E���z�"ʫM!���ō)Tc��]*a��m�.)��!]v�]huj��J�S�<7��=����6���K�����6�n��JR#�}�xT�Y�c�d�kC/m�l��}�A�VHSQ��*��-(Fc��V`���{�G8��`1d$;���%0���;y�m������m誕�_F����?J� ��p�c��y?vq#�-��
��}��db���DM�+�27��A��y���G&�<ؐ0a��4�?���I.�=�<�"���pT�bR���_SZ�֍�
���$�a!��P�c���
H��"r��Fء��\m�_��"U:pp�x0�T�+������y>�������ࠛ�u�運�f#{��Z�fa�s獷J������A��ǌum܁�Vf�tE�'��$��(E�B�;r;����e�u����e����}� �h	^��xx�y�L�~}:>Ju��a��'�x�(�]qFۜ�3_0��0�Gy{C�M]|��� ^#��I A`Y���vU�x��L&v����A�q�-�b��C���*�80A@��	����s�D��u��~'꫘�N�Ԉ̴:���Ph��
<����l���hD���Z�~x��[>��)U��"�{:u %Zzs���ĎL��x�gz{���6��2�,�e)�* �3M���?�n���+��*`m(���'n2�������{_�K-HC
�OuXz�$���޸.�y<Y�֋�e;�~����Gb�$�>Ћ�8�ޞ��= ��M�{X��֢��\�H��I�U���k&���c�#b�n��ݎ��G�~�Y���'�x�	y��e%�id4�qj��N���X�Zh/a���U$��ϣej�l��|�=q�~�;q�}�d�?�!�$������BN�����q�r�4�(={�p�����Y��ޠj/��o�v�B����e�+�p�q�������7ظ�ʥ./J�b�*�U���\�R�K@K*����I������L��?��yJ$2��T�x�s��>��L�]L� 9�H�
0x/���N�r	npmp`&�KQq��"�j�'� �m���LZ�����X�#��%��k�!sM40c�4Pؙ�Y�{S�K��$���u�n���@�����k��;�.��v��}KK^�Vk�92�Pi6����Hx7W����	�BKM^) F1����ߣw�N���	zۯ���}L��ƭ���ed��Jw֘P�[���I*p�^�L��[�7��I��;R@�s��C��+��;7�!�T��#�9?(Y�펧
�(�����?���t�����A�ҕF1�����:�Н+�Y�zIp��+�Q5�+˔�k�E�'C_i��Y� ��D�w��s�$qQYKN������ " �d���o���	�L�����y�y�p!�T����zfܮ��ԮO4��7���w����6fL̍	?�x����䰸��%Q�Ut�f8#�!����7�	�t�hƍ3㖚���m ��0b9>�j�m/�fI�����x�1��Fi�I@��F��&�Q-��!X�[�����lzڶ�zK�Q����,�P	�ˡ�и�7��Xa�ᘘ+�H6"lV9��a]o̞��#to�L_����l\9.������P��[���<���>g��Y$�j)����G\�����Hn��+������;>��つ��^����7Wqa�$���}�m��7$�7�`Te�Ϙ�p)�6�Ε�$w4���Xk��Z��["��p����I�������v������y.�?%��r���!�4��5B�[��!&���#����	J(=:��W��*�9/~�3[�Jע��9z�Ú����/�d��P��$�O���	���D\df�`�]~��)��*l����m2�L�oB�_c��T��|w�߂�]f﹀ ���D�M&hct$���B��ո�+��m$+�=Q6��*�%p���Cg#j6#�S�����P���m�R�X�?�,�r�`~���oW�S�Y��P;�<r����$�tO�܏΃@V�?�L���Bk�Sh�c%��y���;��*#X�55<����ͷbq��	�f��2�԰Q'�n�6:G�@E?� %��7䴉��^�G ��e�S�b "�e�Z���V���YUg��ٖ�ɛ��ʷ����٤�F��fy�Eo�~�i�b�Xa]��i��x�W����X=,��G��_���3:Tt�I�����W�WJ�\P��(;�#|�W^1�H�ȱ�'nY��?��1��N���YҨ���<w� U�?]H����}��(�ϣ-�C����0DH<�>�D.���O���$�pwؔJ���� KPuvW�?���|�G��T��H���F(G�n�Rn@��SBY�?҇[�OC��#?�Z�E]��U77���I���W����Z`�Z<yN��g޹m��"+_5L�Nr�x�v�9�Y"O������7��2hv��@r�u��Q�Z�eb�<����,�ڭ��b�'1��O���ɽ�	h���pLw��J��z6u������+�q%귫�7@q0[g�l+��$���O3��[��]V%��������5f^�Q�?��U"�dxm�b-�/��!�!��)��l������+��$��i����d���w�'~<����dȰ�$���M��(�b�M�ʟ��\���nNK6��ep8��mZP6��(�N�d�@$Uj7
R����L%O�S�E�����9�pctH�(:䳜�2�	��~��m1�a"2�&JOP�l	�,�m`8m���9���P�Y�3 ��F1zR�ףNoh;�"܉_49�����]�];#9�׎Q�ݵO7覴�;���haI���I0�o��xљ��nV��'9�3���1.W-;PNmzt�š>H��3	5���< yB&5�O���C�	Z~İM�(٦o�ƫ�������#��「aL�s��[�7G����o�+[O �3���D�M�4�q-6�5]�LX吾E،��V�\����ôw�dB ��\m��f�-񬯻�7G�*]W��-�+�r���4֤��v��l��9Ү�s�]=�8)�V�f��Y��ǐΚ��	o�W"�A,�n�O�-���DۊҔ�5���զ��N�<���p)�c�Sp�R��x�P<����`J������?ܜ1�iW�[r��/N}<���~�^�B��^��?nķ퍃r��AB#����x�?��_�������ZŶI�O�j�0��T���W�JK���F���1@��K�1VT��Y������$`�����`V����9�f�ڴE�z���_� �l���x灯'���u-��T��`i��j�OOy��&�GX��	���OD�s=�=PB���5�(1��D?	UQ� K�g��	�بk�c͇)\���f7�F�����D� t\�1��]�.���>�Ҷ�ؓM�����������a$��V�Zxh�2�%�=���47�Ȳ�'���c������w޾�Qڝ���z�>�� ��%Ӯ���5ǈ�_�v�Us ���aN���OX{��XnQ�H�D�E�F�I�%\D��i�� �/D�5��3#$7>z��}��e��΀p��W0W���k}v[�9�&�^�+G%��k�`�F�%�����D�ۓ@S	��e��⎎7�e�n�k���*��n%��X�����[U'[�^L�1N.�TT�ސ�)ta-��nF�fIQM]T?w|㿯�D���YS���%�\�<^��$�^��ٖVD���(�>Қ�������P���*I�xPLM�8��j'h6E87d�+BF�}���X�ͬ��{P��0�! �9��b�(�Fb��y]/�z�%-~��X1�&T����DM���|ػ߼%-(|�CAg�1���ն��q�b����4E5�;�Y�д]	T%6��g�ɂ��9�{S���#��Į=� '��ܢ�9Zc�t�)iI����5U)SpTC{H��4W�sTV�V�^]�p�ܾ���UCx�N3�(?��:��ɂ��}�ª?�B�5�h���8`�sW��!��W���A[�bQߛ:6�'�E�g|?ՐSg�/�7h�=��瑘q�Q�b�ٔ�^���}�r���<�6uq5��u��dD����n+MMgd<������ ����\�h2#Ht9xlFM��<���,�N��=a�nO���?|x]��!�݁u��z��y�y�{@���C*6��	����[K~��h��"���Bl��Š�"G�<臸,�H�-Et������Ǭ�w"aa�Ze^����n\l�Y[��)-�My¸Z� �	 y�Ӻ�S���|k~�tZ�:�U"���N܄��HP~�D�$�)
��,�թ/�[5�^f\ȄK�<B:C5�T���X�������rB�/9_��;�<��=����W�G�16���$>n-�,kI;�	:5���{��q:���+pC��?�cbe��wz-���$����@��C���Ub�?�l����a��	�L3���	��{�J�~h��Pz���Q��j���]�x�
%RQ�+���t��~�A��]9�Nrd�~!)�l8�H����:+�z h���]���@N+�a�Rx�E�F��Wy��S�F8�w*Q92btƀȒ��H�V�lb<rd-���B�ѻ�)�l�\w&0B:�W𝔂k����0w����O:��j��^z\p=���[H��Y�z��t}B���o�Z�a�����R~�g��"�Q��@�.�&S��A&��!��[*
4���)~��Iܦ䣤�Ob5�T+��P8��2���Z�d݉��hV,�����/�><�r:H�Րz�ho���G߽��0��ү�.B��� �S�k����t���P������@�-�u��@�^s���k��݄�*\z�++����S��+\U\}�S�meg�)Uy:����g����ʸ�)";�I��%Di��\�o;w� ��� �g��R��xM�@�f��UëG��f1���6v'����L����$'M�MA8��|�D �7x��v�Z�:CF��P}�_�k^�R�bW���F��#���T�!|^�^�5�����p�C�i,:6&|��n�\�*�HI��-�1�tC��oɋ��vNo��5��������b�����E�7Te���ȹ_���D��ĭ\ϫ�h������v��6�2g�Q�v��<]�Wroޥ��Ӣ+����O���QHg���ˇ)ԥ �+9;�y/��&'�A83���+JNZbB~c+��������[�Tg��]`\����N�H$�]5:� `��L�ZN�~iYU���vf����/��k���K����3�8�|i���]�D�����R;�Jɸ+G����<��]�i:Ɯ�� o����k���V{�c��ߣ�}E�SZp�_�Vu��F����i��q�7x���9�%������K��h�1�����:	;Q�z�0�mGN��D�`֋������8x�{T>3��K1��i$qʑVN�y����nG�.���ᜂ�(x'�� ����`"DzND׶
e,�kK{��:x�Q0H�1�3S��Y/M7$�_J`�,K � #y��>π�E�3RD�nq����`�X$�]����sizO�%ۦ� ���b&��8{��&]4)�a� �da�HL��k�������vpG���~`&��-�f�Ҋp�}6���8�lf���d�R��MJ�վ��`a�4�G36��-�e�WwP�~�a����h�8��H��t�����/�r�6��@h���f�>P^�;�B�)�1��e�2������j <x�'C�I�i��s�ڦ
�MŅY��'�ꚖcOqL��m4%`�{�q��^]�{{6�O��U��U�>�����5q����i?�9��b���]/f��e�n3H;)�d��"�\9r��~���Ks.i	�g8�����
�6��],�h�_����	<��H{}��Ն��������P)G}E�4/H���'��a����&98̹��`��o4`{��ͫu��A�{ɸ0ty�X�K�	�'�|�;Tpa�_���K|�ꃵ�����X>��g���Y8Q
�YP�푈�"o�C��� ��=W6Ɨ��PW<�8��衿��)0�A���v�E<s�9�,�6 :���1F8�<�A��_�ʥ��$ \�8A����Mʑ�'V��7�d��D�F�x!1�L�f^Čn�c^9�$�H3�� I0�+� *U 	���}&<� �m��;��t�w�coLgPH�`M;7�`���#��{>&�+ڢoR]D��i���F1S8Vl`+����|��UR��R�_�iNx����K��+�e��z�FCf�ծ�8y?4sqe��Ӥ�,�WG~
���;I�x�L��$�5X�پ����M��ZR]�:���o�]�s�'��&6�g���3P_U��F�t��K���NE��d�����e�T�:q��tű�v�Ț���Yc�E�N���h�!��C�����?�0��#�*�ȽF��Υ��ԁX���E��v�nݸ�ƙ|����"�r�8�G�;����.����d�AWb[N�M~%�0������%l>3Aθy{? �:�^kQ��"�A���x��ͣOI�v��<X�E�/���X�Y���Ӡ�u�6�o}k5S��z5�i���gZh�'�~SS���ؐ�1�>�t�8;�$ЧN�P3���~�">�>-���$\�C��Ǌ7LpX,b��bVٳ�,m(� ��W�l]��IF�p� Q���%ǖ����άy�z��_&�sy�p�\*nh!R-`���Kˌl�vqǚ����M��X�5ʬ�$����n���O����������H�j�;��Z��s��8K@&�s>�����3�?�t��.��Ar�~`�����ɚ���d$���t��ۡ&�4�in����V��AC��N��H�je�����"9���1�(����2T��r2��� &����Sg'�C`r�~s�Y"$�����S3
h�R賏BF��+����� �+R+�6�N�wm��>6�-�$�t��|װ�~I/V�Sї���i�ҿ<���|������\ː�P�����]�:�ᴦYN-:�'P,-���a}�%\����_�[���]I&!��#ߧ��)��W+�A~G�-�
��Db���(�t&�4U��+m��>Z��֡�́2>L;�,�FvK˻j�5Q�e�W�&@�A��"4�
{ c��kG�>ŀB�q�����J�2������o�R�%�ޡ���/�=.�i�JKH1� `7�`B`ш��*��1M�y������i�o8�ۘl���g���9P�ڑd)����G��u��#Q���1Q�V�i��q杏��Lk��Ğ�����27�%mw��1P�@캓�Dp�r��{�&\���D��*c��۟M�<�`*l���e��㰢�G��s	��+m[���ޢQ������Ug/VBWn�I}-�@�t0�� H$c��3�}Pޞ���x;�z���]�ҁ���t����%"�џ�rD��Ø��K�>�����zwl�� ������	��t͛�4� $a�j����Z!���W#�u#�DS�F��`�}Ն?�Wsܦ*�,�j����G�~�P���T�9��gM����%-F?��^}��|�'Z�����C��p���66/���X�#���1�.�d�w����a(~/"o�JXY߿�mp`�댚���t��[���~�ا+��,#u�F��Y��=|�Y�&��B��"��vL��5�!K�ˈ*�Rx��a�*�,7B�kR�"K�2�1���(����D<UP.ũ|+YAǞ����!Y���)d6ܘaR������+���n�������6L�k����E���gX�*��HN��̏p1��x˩֧c{�52eE~��E�um�M���\�� �ڳS�m�2�����
{Pt�����u����O����v����(Z Mk�.y�x�ْ������e\���"b�l$�,X�����x QeS�[z�k�Ik�s1�N7�m-Fk�aD�&=|��,]MD���l[���q��yQ���>��b+��c��$B7L�Qϙa���S�*Nx�~vt0zj��� m�Wٔ����$�@���6E��MU$f�~;܎Y3v�������(�}�\���^��ݨg���+�Qz4#����o���s��O��m��yS|k��)�D*� ���Q{K�;q�=���,��N��KM�<��7*�\�
�HlR�A �E��]�7����� ��r!zAE�.&zMϔ!f����	�ίZa���C��^vX�<���F3��9��Xq+䈑*=�OE�v�)�u8�]�L�擃=!m3O�r"�#}UV��چ!�����>k��5��ċ�����R�C����(�؋��l�/E�~�נW��=d�e��ss�ٛ���r�ɟ ����`2s�"Ku�z���Hy����[��N�}�lh����u��L�{���5�O\N�U�INw|����Z`=��,����9�g3���8�.��>�?��M���Gj�ѭϮ�Hȝ�2K�����5O�l~_�">�y��b�hU��E����
��@G0i[��)7����y��ų��&���18m���cT�l~�Rɇ�ڃN�ٰJ��a  �~|�b�����	_!j��n��0e�.�Nw�$��u?�n�!����䞷�_q�<�984V��������%��Q�w�G�
y��mYԓ���@���E,��I�)�����ި��**�ݝ��J�`������e�B� Y9�8��,~ ��jL���{9���z���"�Y��;�U�d'�~~r]�	]�w�xg����\}���:j{���f�mX0�B�s��$��`��  ���#71;V�W�k����.INc��3K�y�y�'Th���#"��ք+}�x���G�?jXO5F4�L��1����h:<2p<IY.
a�Df]�U���D���#���+ȹ]I� ��g�<]MM!��] F+��ۮ�Ѿ�b�L����+%G��_��I��p#t�r8r;Eq�l�i�zo�J�;�_���b�T���H��e���e�<ܱ��G��K���h
z����Td�~;��nm,6�d�߯�!�I��%���_�$���~�t;'�s�Zi��g�<4�sI�}�T�x���3�I4��3��"�8�)�4tpV`��`"g��D�1��2wc�|������6}�(�u�5�k���PD6��b���t�c�W�k*���C������1.ܸ��`@�	���`V��0;d�g���2�����oiuVn^FAo��x&�'O`R��1ޟD�fh;����-ř �0 /��`����שˇ�χl�*f@����9�B��D�,7�����y<tC�	KL���.q@Z2oޭwů�-���#	s����+���#c�����7`P��n1Ǽ���%�Qv˒,c)�����E|J����]�Y��($�vͺ'���(Be�3̭pzb��&����\����p 3�ca�EQ�YV�͟$a���,���/JNғ����e#Z���RtTo�耛a�rV_9hu�K>m��ZGB�P�Ofַ��x�1�!���G�Joc�f]�μe"����V���lG��yAbaD3���Mh8�eu ��t/���Zt��
5����6������*x�*O �h����7P�t~�#���9ўk�*T�ҫ�q�=2n����R���P^<��
?�^�1�.i��t�V�v._`�@ffJ4W��(��N��\)��2���k��pt~���ꈄW�kv�,�l ���i����[,c7&Kt!���X��F�v��Y; &!���5��ne
�~{Mܯ3|{������Є�g܀���p��\b *�@����� z��n$rE���d��I�U����
�y�*����	>Nv�N��0Lw��(g|�Ẋ��k�J��<��sp���C��"ɔ�͕��p8/��d@�$[��f��d���oq��R�}��h��$�w�j�i�|mq-�fӘϻ�vƺ����/�����᭩:����EDelǈ���»%� Du��r�����ƻ��4�p��M�F�$��$P����&6�W��3~��H̚<�3��0�M$k�h��]��V�US�+޴(�8�h����m���@���K�5u<J?�2n�Q�Y��ѽ��DG)9Nӆ:���jmS�43��)/j"�&)�M�SL��Yp}ůJX�/9/�3Q�x��۸w`I������U�N��㽺f�����+��h�{�j8�Ńf��1�٦� ��n�͓r�����3��B�O�v:@�����^����8�����?�V�Sfg�3��t�?����O"�Z5�T��u�,T�#���U��K3� ���;|"����J���X�>���j��Bس�ee����^yK��m��	fl�ׂ�_���޵uvQ*�m��~�5{�q�帏P���H0z�B�.��[�y�������U�o�ȾR�w�pe6�.:��[�O	�>&_W��K���K�b*�� ~�>���A{�
�c��gmE ��_��u-��O'�'w �X����b����_��-��H#� %PKl�{��r�v�l�����'�K���5�L"(S� ���"�p1�`ʨ�_�;~:
�U���d�[�ēN�m姝�zC�j���DT��,���$���҂'�c[~C�3�[�Q��P�f�z�^�!�T���`�XO+��<�Y-Ԧ(����^bh	5O�f��9� �����)s�X�Ba�ǋ�����|�l*Ej؁�$4bl�/v�1����5������i��7ydCz5(�t�#}4�v����ߤz�k(�� .%�K�ȧ`�!�1Ժ��_x�j�ܩg����u���Gq��CXeO�{hje��8�)[b�7�Z����n����gN9�t{V�l,6`��;��s�w��G�S]����g�{~j����yQ;�gh2�:�' ��]+��шc#% P
��[���43��WЕ���k��K�^���>���#P�ۥ�7r��)r8w�����9��.�J_�>LR�	BWt�G��{td@;�My�Y��EE��N^�xIBޫ��GG�(��At�_��"�Pb�v(q�3�{O��H_"�7�2n�~`9w�ب\��t��v�y�����̖qj�����$~�憜 ]/���"`�b(zi��sU�*?����D��
N�����d�:QӸ�a)D�
eϝ�ћ��ǠJ��NJc�cW��;G���,�lND,�)ΕDP�� ^�p��&���x��y��
�%��ٚQǏΧ=���M���
]U����u�Y{gn�2��7k�r�S뇣�Fz�\ 9�p�E7)a&�]��:d���u�Y/�p�jaq�@�<Z C%�6�<���𞢠��#r�����R]B������ο�<t��T!	�K�/�=�F۽ok�4��kT���u��T�Yo��ZֶR������1�_g����!q\�`��.�R$�ؑ�݆-���*�`�p�?޼�}�.BC�y��<�CC�-��|����$ue�j)jy"#��H�&�����c
A��]/��  Q�g"�6�}��t�G�r�{�R�i��4�������XN��s���yv'���@�F���r�$1g� �堎�������|J�f��i��z� =h�qd4�E����R��=��'��7��t�	Mk��{"�Y���(��wC�䊽�9�1���O����GI&�n*��4W� ����Yڮ $~&�F ��Q�e"��D��}�w����oD�>�^z�pn��Z9�M���ŷ�r�������~��8�9��Z֜��=�Me��a��h� �:PfF�B�w*��_�W�Y�˴�'+H_ 
��*��"7Us��e�n>H6�hv8�� z�wu��Yä��Z�B��G���Yh	-(w�����H5bGSp��{'��FQY
���zҀ�X��5��zA�ׁ
Vn�1��$���M:��͛bw4E��8���	�ӂ��#r����p��M���9gA�_҄��o�^|�����B{G�-hV�AC[�u�v�q��H��y������ʌ�mՠBk�L5��2��"���FG��c;nfItry�G��4&ѫ����2�P�ĭ�`�H�Y�C%�H)����x��<�'T�KU-Gl��~bs�M�@]ې�Zi��gch��-�.A����7��̎��.����ƜD�%���_?��������Y���O�u鷛U��~Uy���������k9��b,I�b��k'� ,��@cZ]�Y���pƚ,{�hYc$�@MLY���{E�V�|�ז����a�b�G�=��C���XF�i���x�G�p{�������1%Ѿ� M�g�\7/.g�`�c[�	@ȡ��L���;��:+�����	<
>ݚ@���(>��Nǁ;���}���]*��j��&���Ȅ�8U��0��W�j�kg1m�L��%T;�:-p�(|�}���B�ύ2�t�>���M�[ I�cQ���+�j7����.�ʴQ��k���6�(r�7� ǹhSr�Kn`ū��C�~Ծy� �A��=�`E��
���T���
�t��b�l�s�QcgY P������\���_-��=��]5{18����hɯݔi0H-�=�ܚ�kw���;����D���=��+��Y���@S�EG��F"U�M"M�>V����[i��C뱝z����N�
�1�"v�^�G�q��3sl����;���^@��9B��*@��J�����nӸ��x)?���~j�?��l���m�?t�g��Q�Iv���^?9T �i����­�6�^�iR�v�[�n��%��d�becB����ߡ����M��\��wK0Ϟ����Y���Qѩ̵i�3&��6ْ����_�p�N�8��6��B��6����9���P�b0��x�Q���U8�������șٓ�/�ɰ)]�؊�G���p<��T���0R:����.N@r��ӡ߶��,wq�M�5��!]�OM�㙢�e(��� N��U���~w��@j�D��8&1���V���|�V�ˢˣ�_H-�_Ð��t�a.ʼ.�q~���7�����*�U���M4�yd��c�%�c��Q�����
�i,���Y�5<����]��y�T�Es!��	V�V �[�3���}�AAoQ�5���U�������6�� �`ۅ��zȯ}�y�_�$����:��1�����Ƅ�n�0�"�,�jЉ��L�GC�8l���!��)A��b;F�Qx࠶/�'�
z��:$:7�3w���$A�����Ih(63!M���᱗''=<�$�)����D�asT����oZ��jy��<����&_߉���o�&��L��҉��<U��[�#�������h/W��S�%�W�c��;t�9��G�S����۽���FK�$�y��3~�Oս������r}D�{Q���W�����WY�wRY�;�����R%x�`�+�HR�a� �]5Gc�W\M.LO.�|K�[�ƍ�)\u���d��������ʗ�o�eV��r�1�XɄ���%��ip
�3h�p?����f��j
��A�S2�._v��%���.�k+�jfE��Yo���de&g��M����&3n�KvR]� �Sx)߮v��(@�A:�d��.m� zkJ�du%m�)��8��]���9�A�S��l]s�[�9����Li�(XAs�5R��y9zط2�'�5$-�ǋ� 3l@;jQP��И��� ��+gOZ����F`�d��݆z	���p�$bN9�&�w�#� m�5j�z0\Rz_���N�k@���<���C[���T�`!�\l�����=�cv���y¬m�n����o�ؖ��,�bxGGi���NFwr��U�"�vߟHBVx�8��}�@,�:�-:�`�8"��r,)�=!j���[�����I4Jۡ�e��{���+찱x��}$�T���C��(_��ǫ�#W�$�ދ>�������6�	Z��qބ־	�O���b`����S8i�q�����,yZ1r��\D�����z�CP��4�i��P0��v�`�SY#0�A�-��s������O,|l�/A���~�T}ܮ*�D�~�"_5%Z��l���z g�1MIA+�jt����@��2�J�[W9W���5pE�׬�ʘA�Y�]���/Ě+���ȝ�Y)5^'���Sօ0ճ?:;�P����RvLԟ���4�}�O��>��������Е�+�ѸP���F
Lo.PT�CR��'�"����q�F#b1T��3VM�3 IoJ��ʅ�J���5u��@�gD�/��� L��P�a��m�����ůa�L9̉����Y�P�s�Q�G���n�@D�d�����`7����ra<��������mă���҃Rb/�TFȜ��֛y� pR��s� �hⷘ��e�?+9DU����c��T����R����܋��d���9�,i%�����*��o~�CԞ#���#������'������:lþ�1� ��Kx�����'R�����9�
��J3�ګ�o���K�0� ������󪗌S�Qa�@C�J�a���C�����}˷[Y��}�B�@�f[������V�\G��5���u����!N�R��c�:�n@�
h$\/��E�,��G5aI�c�G&�g���𓸚���1ک���w�ݷjƗ3����h��w�:�
L��<\�� ��4��0VϦ1ұ�]�w�g`��0G�Xx��p�,}�e+zJK,�B��UM�{Ӷ5gG��	��� ���������%��eM�p��
|s?�����=ֆ X�Kkצ��滺����ߕ�SwJ��K�}�RCt'<$T �);ؓ��#�3�i�B�_�+ o+B�"�o�b�r.R!b���Lj-���u�~E���,W���`�ow�?�1\ �Q	�B���u:�����j*H��Nzzp)��1�r ����\�@G��r�:
u"������ai�+��f�=,��x�U�>r@-a�IX�+Bǐg��:^e꠻��;?N]U'�_���鰕{b�Z)u�w¿G  r�u�l��%z	��)�a����ה�xu�D�(^�����/G[[�x3���p�;z ���D�0n4@g #�M�2���[3CHS�?��w �Jo���2�}����]�J�ZG��X�!��g�x���Vˡc&uJ0����;�2R�qM|�qW8�jzf�&�C���#)���@�=W�m��(6�7�#(�QG�PO�C5��a��`�nV� �Z��r��晬w���I�
�9�v
�����L���lS�"���ֽ-��3�q�O�O`�����gRw�N`�Z4��T.��A�L^1'�R���-+p������;�I� �781�C����ר����
��ƲF�e�+��,��>�.��-�0q9�dٕE�Lb/&�N���{	�C?�/5��Ƃ7р������j�,5%
��ʟ��b��^�0EF=h\Q��ܥ�WlƜߡ:�T}1�~m��� �}	���"�V�Dĉ�U�I#�5>_�ײ
�Zߧ��a6�/l��5x��[���ܯs ��	���b�����:�?��ne���"��a�T�5R`^���a����Y���; ׻������#�O�eL;3.ӑ!��� 8�'Y��  ��{;�5n�ܹ� *cd���D|�$s�>��:��y��0�׺�� ��O�a�B��}�I���7ƌM%�f#�.�E��i�6x3a0�XE���kpF��m���I*lB��S�\Nq����n�����X_�ev,�
�A ��3!��\��$��m�F��h�����譟��[���Y�~0�v�w�!�Z��R�Z�|a�1Dߔػc��-��ז�9�-���{-�03~��6m ��,���LKC�j��c�}����Y���xF@ȷ֘�(�-��i�3���^o�����I� ��K� K��gE����`��#��j�l���<D(�9�_��g��)�z$u���"�r�TPD�^��=lP��Rf������H>��	�)�N�\O�.Aa֓;�<�W;��a����zVmj�;�q�Z�vv�����
���
��4zJ� �2���3�ř�RUe��%vǪa�9�.�$��$N���濔�d&{!6N�Zpia�wEwѝ.���k �����1�����|�K�X �B��ۋo�$��,�S�Q�W�0)�8X��{s��i���
2Lu�3^�`�f�� ��P %�
}T4�1G�R?L���b0ד�/�j�"�H�� *���AF�լ�ad� �i0�O�y]�6�x�EB��R�
���K-+�*��|1��V�h��fY�?�<P��R������Ya���P�]��Jt4yo�M*�CEt�E��x��lRT�ҏ��::�d%.!�~�0͊a#�|�N�	xX9S�n-�F��KB�7YBX�2�>C\�T	�J�L�Ǟ��<�kV�A�C�w�6�*9�Q�({k�|F�i�u=@�V��z��W-�%{����T��
h:xIX^wC�g5��x=nʡ/a��}z���j��-�����@$�1��v�-���ls"=�1�@&3�'���Q��h��Ok�WKƼ��]�9��sB�z+-R|�Ӓ�6��Pm�`���EA�P6x��|�z�՗�"A�C�B�W�a��/`�H8-aՈ�Ν����������KKKfl@d��EAd8w�l���p���;6��ZK%�T���^0�\p.���T�飘�d��6NkL ����RT�(E��9Q�����9q	n��=v��$�@��,�	>�\^���J�]Z������([�w������0�	�o���f�B��1ǥ.z�:SnSS�ҍ�"ŧA%B�ʎ�O�����p�U�f!w�T��vk����^��J�*�	l1@ԑUv7�|��j�1�O��׀Go�IN�Ai���@M�ޜ�����\ɹ�PG�~�ȟT� {^�>1������߲{=8n	T�=�mʟ��.2/�/�:����-����S���S2"־�MXm
#Vc�v̘���
i��~˳���#�v��f
v3��`Ȱ��y�4�r�M�L��f��:$	�;��i��"	�u�>��*l�S�KK�R:s��M�T"�U�G̞���ŢS_>A/ǷsU�em/a��Tv��+�wi4D��j��S��_?�d뉉}8)��T�3[������*��g�-W�,y�C�RJ��s�j���r��Z����CNz�fV6|�{���`��*�{yX�����H\l"���v������i9&g���LB�_��n���]�$���Q���k��C����y��(�H��7��x[��@��np�e#hX���E�;�R�˪�9'b �N(���W@���B�H�P&D���	M����ˊ�6�>]F�(w��f]y`E�����O]i��q���`�8��1��F*�n�[<�9��y+�r�� 8�N����ȭ4���/����gN��Ԓp0��ة#�6&|���lqts0��P>bW��	��x5��agTN���r)EC�C�������~���3���ݜ�ʾ��L��o:�Ui����m;<�Q�
!��}�^ѥ�IeY��E�ӲI̞N��i��bo�F�:ur���҃	�b�Z�@���7h�]�LL�k�	r|�m�`A-�F}�a��0e{wI������H��� ���
U���Gؕ��H�Z	Dx����gw�c�m�'��ϊ5�z��P��K<,�<Al��dr����@����$�#��3�\��c+�fmf�����V�_����186uS��a��� ���]���0%~sQ?7�	��k�=x�oV�B�n�����e��9Y��~.?�E;�g
�?�=j�+���p����yb���;#�xf�^"�ڏ�dr�
�����s��-m�>���X��0�1�$cݟ�3*{�&��>�_�8 ���U�u���[��KC�΁x���4�'1�D;FX��
���Q͘(� &@&~͜��Ak��՚�8� �N ��ѡ�g]��c�/<�r�^/��ļn�]�a�DZCh��1]a$�\zI�͆?�P�&M ��o����"�����G�f�Ku���k$*��x���m�O���)�+`�TB�����|&�ӊ{f����.�Ұ��M�עa�Z�·�����\k�x4�y�('��E��eB��ڙ��=���񟖸�S�L��h�����&lIi
�z�Ȥ�F#4�A�����?�Һt�h� �)-?����?�I���7�%��O}�I$�x=�^�H{Ւ��QD�nB�f(��V��J��t��m���o%�}5δ�<<��l���yu�Ϋ<8�,c.`��&I���@�x6�{�����@Y�e�$�pTA6|l_*e�$���ۣ%�P�o�S���-���t?j(7l�hK8�����>������cY|�M-7�	��I�&�h�2` 㖲*m-ت�����vf I�z��U]%���s�Hd�Oj`W��e� �j��Ճ���@&)�� m��H���$K�qY>#;�:�c����ʫ��\�E�rS=��\�̦b�4l���
�K���͚Ɲꗦ�L��0��D�.g�*��3K0�w��Cd��ZL��~�Eiӝ�߇��� ��;h���W+su��5�7E�o85v9��,IM�8P����P�+��8�?o����V�5}w�L1��c oJ�
U�5v�f(U�����B:�*l�J`�G����8���	��?�8�Y�k�W-&˸;FZ��4�g���H���{Ĉ80-�'r�����ߪ1{���r[���ʐ���-Jg*&��s�Ϭ�&���p�~~{z�3�+_+v�C��C����-ڿ֮J3��lF���4�Kjj���#`��
�T�,_��\U��Aի�͚@�颎�-�x]��{>�U5��*4#�Z"#�0��2�/Ɲ��Α�#{� �����-卦���l,��P_���*<m�O��ꄩ˸���?`�1��_6�|���B^��vK�텔��RO��v3�n�!��e�B�Dl.�ew^���%�S7�Yn5��ke��1<�T��^�o�禮
l�EJ4��*�U�;~�uC�}�������$��m���wp#�!
�����UV����|�!�j#���s2����l&�H&�g��2���F�����\a����WT�e.SB p����s#�DKٜ�$^�$"e�<bG��夨��ɸ�X��C���8\ЍjI�|0�Hu�|�,g7� ?�D��;���ȐUb{�z����0���>$t�q���`���)Uu��4����2I�ږ�W.oG��U���>�!��^rD���C&*�0�d��� )R�N�?��;������<aM�9��oF\,,�s�����4S��{%��\n����=T��; ����c4cv$�& y3Pa�c��9D���\@����4C��.2S;�'_� (b�W+�G���}�H�2����wN����z�_�3�S�:��cޱ����Htk%e[&��0��^�F]��mRQ�q�� ��o�����%,�sˑ@��ЌQP��}�ޞ�H�ÅaPa��ɢ��.pWFsH�o��S���v�f�f%�k�o��$k��-=`��������A�]�L������ ���7ʗ����(Lc[�붑�E��`�"��[.��m���G��W��oY6��G�m�D\x�(U����k��WA�����N�JPw+�n���=�)7�.d�<�����+��w�DG-����>��Cv�T`���5��a�Nȵ�P��(kI��I� �P%�7.B�M� @V�taC�ˑ���v3΋Z�
T�tn�Hb�Ж��w�=��r�o�C�{���KW;6o=r�8C�sS��2�3��Q����oY=]�Z��&�������ܞ�c �P�������N�������(�c�$�܏!�D�c���еRk&��p�A!e&��#�H�e��<�������g6���A��TE-�X��-���]�lH^�Ql��\w��]��:�{���e��_�
� 4�%.A!AJ<Wvj�"ɉHghvN��;�1�f	I��}�G���;Pk?�~Y�.W�#�!����4�UGՁ�K&yj0wퟁ>|H�%K#%:JjQ(�Ԑ��#��D�"�� I(�G�l��hW���"����2��������b��O�
K�_n��!Vt&D�T����$�n/�m�tXWT%�y�(��Cb�6`G�2|��2�2��kV֯�תҬ%��!�����+�*鄆�]�w�
��4�e��o���w/�����Q��/��p�n�9�r0�r~^���/��m|��2�Ӹ�]*x"9��ș����A����������F�x���;�h<�:�Y���6��r�Cx8}_��۝���A!���V^�Vj���ι߶u��.j0Lh��Vp��E��*]�5�!T��
+�(y�K�H����!�t���c���F�n�}3/����c�/tDy	ز���E߫M�U�@C0�/7?�Tf�l)����?��e]����l�^�V��������B]S>�f�j/4#=V���<4 #$��	�_l�Ft��M��~L݊��X��[PE�?)�!�²�]F\t���9v�@	��Te��sd�c�g�]���_A�&�Q��i����;����`qӤ
;�k��#�I�����4���)!�ʅ�XLz��1�_\���
�+v����-�g#=�vf��6��Y�`7��6�n/���y���� ��W���rK��ku�v#m�}t}���`�V�Ճ���!�����Qǹ���V���%�UɊ�SՁE�lo�#��g��s�
}Bz�:l�%�~Zh���'�tI*���~��z5���)��$%��M/�̵�
���;�����)o��/7�$�92����=�q�iA)�;�%�V]BՆv�M-�O]V�|ʯ^�NX4�����+$?��f�R1!�;SrV0�0~Kj�W����u��D����5����Mq��
�^ld��J���Ue��`�l��g� ����+�\�
(��O|9�$��x��6�#�V�L�4pb+
����(��7h���s�( �ǵ���(�_
)�.�
٭��<V�#S�n�5�/]ڔ�����eq@z��{'�g݋��T~�W���"��kS(���� �ݩ�'!�;/k8�?gK�E�]��5�Ə���+� WfNLG���!�PFZ#�g��\�F.������K@��D%���.ܙ=�6@&���ڶ�DD�i�]:�YKJT�n�0烢����U�	��; �܈�(�(����_]@��K�{�Uu&�y�@,��J�yi:t�>;�!���Q�M���!���`���4�&���e��I�z��.��S�\{ib�E�<(��P�7Q}�����j�����]��5��<��,�O�|n9�u�g�`J?i��5�D~��&�� q�y[���\T��q�E�謥,ؐ��dBI-awm���S�Ds�c)���P���6&��X�ݺToi�K�Q��,"�z��I9��X~�<�i}��c�ϲ(ÿ-=���@}���I�e=����H�"��|�n���Z��%�VEۢ6�es�Y���_�r:d��ݣR��hR���l��}�v߄�p��$S1/'�G�4iE�s�%�t���f�#ABd��\�l����X���&	�*~�*�b��E�z�y[��L{�2#2�HFTWh+����+�󬃩f�bϤy�l �i,��~WK �4��e�#=��f	��3	�0-n=ೈ�����:�>wIپ��7�Aң�8��|�=�b/��jK��3p{.E����j����ge��@C� �z[�-�b�O	�E��<�-J$%�*��
���E%�|;E��k:��e@�@D,S:|��J\���)�]���A�4ǈWJO��$�J]7���t���䏉��z�E�����s�Ko�<ū�.L�?��&y�%��}K{�#LFȁq4&N��yNtI�9��V���k�F �f���Gjˆ-G���3{��x�Xg�[&��&k-y	���F�+-��^��2Ci�Dš̞܀��7�C}�~T��.8\s��Y������$����kҳ���y���q�}`��ڀ��"t���%����X�"zb�c�܃�e�F�H�x،q���n�y�W�)Ca(� k,�h�����㦀�Y?��]S阹IM��YV��W0@�e@�/n´�Z��c���e�:��Ϟ"5�>��~��o�B�j�H�s�����'���$L$�uPZiAߕ��@}����b/�s��]L�yt􊁯��h�k��a5tb��z��j��4�nCQ6p�N�(�c]߼j�8Ir��he��L����˴vp�0���8s.�(�M���ͧbG���tg��W{��w/���'ʺ��M�ED���Г�Xpק.ƈ�]::r��<)�7T0�'�1�넟g9k�@*�����O݄�8�����Ge��}�v?�x2��0�K��xG��M_hL���y�
��p�Ǥ8�L�jj\�%^O���0�~`u��P͓��ǝ��"�9U�,��W�t�T�,��Һ]5�UZ����Xk�YiR�U��:��i�}��#Y�:�}(]M`��풭��,�q������L���R��O �l+��q�}������:�Y�T�jmA��m��F��t�?c��Iϙ��qCvZyzx���)\E[ٰ�ƾM�KyN�N�5$*ގ�2��τ��St����CT���
�lg�	��`+#t{߷�od�jF����G��#��E�oz�&�<������Z7{t]-�-�#��z[˥��$�C���T�?t�#�l�]% 
��"V����!+�|n�x��mxI*�� �k�bb\���q���>�1s���,���DE�����&�L1���'7(| ��nY��+��&$'p���hx|�8�m�F����9Ȣ��#�b.�W.Gٴ��I���^9_?������/�}���9�����,y�mO
�P?�b��|[.^<�,0��7 �U�v%t�]D%�)�ȤH�L[��i<R��:,d��w�y�e9�h�,��c���B[׽�0����	�II	�}�uF�6�$���|���k�0V�D�PЃ�^�l�b�#<*�C���>��m����U����){�S��+��6���?���8��Ca|��q(���ňs���Z����Uk��^��j��R���k��b��zV'�Gc�N�L��X1+�X�Y������g��Hps�wV3����O5� ��$��:��q]���#n9�ehM������4Lk`}�(^�#ҙ0St&sX����3M=����pK>] �7
y6eXB�f}���-���cF�	Fݛ�l���\9��o�R���3�4Q �v��B�q+��;�a�N#X	2���V����kv%�f�S�ݏgf?�es&��7\���3������9"��dv#�*���wMD��(\ߦ�n=��-^X�ko�;c5�ב\��e�X��:q�`b=���rL�I��d�oO�:(i.;w[<����<.
ǂ�#��"�:F�nܦi~�v�b_3��A�*��c��^	��r>>?z�A$r?kҎ!^���Wk�Wds�h�D^ӿ~�*��܍D(�����W�`��Q�/ԼFڐ�M�E�6�ؙ���2h��|�KD�%�)1ٛ�y��%���&��4*��# �Ē7��rJZ�s�+!�|܎ ,�N�ާ��.lSSx�$���eD4���x���	q"�A|w��\N�q����	z�V����ݴ����@*�FV�D�EG�n{�J>FD��'T��G�����e�1�<��O �@�qw�7ۚ�
�9�Z®� 4��O�.��n�Q��އså�ڎ��8!AE�i�˰���=�'z>Ɣ�8��z����`��S<����O�7K�I�D�K8P�i룼?Y{>apf{e0=17+Z�3�R��m����ɳ�:��3$@��潩=�xRT��$�s(D�HLz����YQq���⫄����<�� ��7>|� C7s��t���*�ʕ��ө({Â� �5u�d�\�����FN��~2�]Ѷw�C�J��o5��Hgئ�g�!�~ƨW��[55����d�:�iŸ:�/�R��㆛<���+T:4�&���~x]oi�����w]#�҃�^�P���b�h�$�x�Y��W2 ~���]�O�RC}�|�k5P�"�	 l�
�<�S!c*�����#�Ʉ����C�H`�ю���^�XX�;�.�$����K�k"���L�Й�+�X�n���a�؝㷮���2b��iE��.������k��i�x��ǫ��'џZ;��ŷ[A������G����%�JGI�;���/� !do^u����\(GG�~���c���$�1VGd8R+�reÕ��j��6��9
Fq��
��4It�%�Sz1��6����$~��:���}���?��P0�P��f Qx"�Ҳ��i_���D&�����kq̓=`�)�4�YOD0F���"н�?�(\|}�u�"�<�W}B*f�ΫG5$���4bKU]���h��<��\5&�w!V��H^ VFi*}��f�AdkbN]Jv��{�����p�8�4� Bx_�u�J�,;I��M�Wu\�D:*��bmi�y� ����R~nb� :U�#]�		H\1�XNg�2=FBw�X�Wnm�Z�1�|���h/r�%�al���ߕ'!s���`'tQ:��(W)��w�yJk�u��>�QTфr�����y}��|��J�����N�i��nu��R4_bkDp&�_x�LvF�m�7�x%Oٛ�Z�2��PgeK������e��{�R��gÁ>!T��N�8�.ŧa�61�$c�l�����M�wm� �}l�`���~�Q ���_[��f��PK�W��8�q�j����XkG����mZ�v-&+�\��]�p� RT`�xzw,�pe��ᕸ�r���#�4ܒ�&7�{���*1ښ�v{RW����ڝT!%�܉�jQ���!L��갩^'�.�,�~�,��������?=�y/�H����9��H���Pi�Wn'���!�֓�y�X�
���\�ݼ�J34����7N�BH��R�H�����W�0 ��ctGǢ�[�� `=N���4��d�M@�l�&�� ���v--�)}>��и4)P����_��#�/��_R�%��!`l��p*7#O��͐�[��hߌ�+M�{����+���f�@�V�8.�l���{�S�=S���/~2�8@0ۄ:��b6ZX�� MK�X�|g>����V��s�+�N��E�s�,�7y�%}	���c����j����;�ځ�;��;mpR���/�.M9����י�kĮ�ī�|���Uۅ���͜�+�3�����.�^�ko?�:&[C�M�[�U�0Y��g4א��q��RY��"B���g�_�����������r,���q�t#o�<W^G�R X"�O�'�)oS#8j� �%���sR����V�M9�l(G;D��}�5Nz�l������nݽ�I�`�MP^��`�3�gs��ʕ���ϴ����J���dpP$BH1֭��ߕ� G��-���l��7 Aa��b�@P�k�_=��%&ߝq<.���k��W|Rk.rj����PtpÎ���G��� ��&��ɩ������ R ��EEi�Z%�����#+��Q�/r���|qq��3����o<��.���K.���ȍc��l{���6{���z�5��q�[�� �^x�TF� ��8XZ�B3��;�bEF��.�˶����p�ރ����Z�
�s��\'y�q9��f�������1*�w'�&aw����̋��3]��w���߹� ����H(Fc"��1��Ih�Yr�=�ÑMD���&�\=�`�p����|t�GӢ��`-.�̜�NL}q�FQϝ���Qk6���?o^Մ=n37C3~j�7�?fY
������9����?&����0�ib\k'��ὒ5�K��;`;G�
���P<��r[��Q*����+�p�%d�����^P5�K�@����(�f����UV�R���A�#��01��I�v�>��xl>{������3�z�-��L�EkD����UX��p��l�7'������u����]a*�;��xl��!_�S�Z����^�4_�����ꤊL��(\�ۗw��1�Z�1z	�Ia}�VM�4s��Q��0���C
��ߌ k8]j$즱����z�lc������#������1L�s1s�8e�׮w�Wz��%-�opdOS�{�����&q����_�c�?3Z%q��\$����\It��\c˄���Y{~jV�T�	2��@�r�hrT��G��eH'��Bս�&�n]Zh�<�� ���Xh;�/$%q�1�q	�$�ڹN�$�Jѐ�1W�q'%AL0��s���A���O��������R�"�F׻̺.��`Q�����i�o�$$F"���%�`q&�Y �c�^&5`�0�SX��D��9o�G���&ٻw�g��M1(F�LPjNʭ֎�>��.ǌ_�w�>��'��^�9Q*!����죑� �9�п�`�f]̦�h��{5}4�jT�@��sS zI����@[U�[�~���|=^z�[B�+�J�톈hqXUI��0��S� ���t���A�K�2�`#
����^���x�*��Rl�(.��[4�OD��zl+���{BG���+EO�Pɺ0�I-���f)�΂� �b0��Y�%0�(������h�W���!��7�=B�B�F�� ���
[&�uy'#1���Z��oh�Y�4��eM�sq偍1/(c�k���Ыw��L��n��M�9
���Z.�nz�u��8D�N$9�x���0�I̺��lC��_�+W�_�Y��q� �ue0��ɣ�2��QG,����X��6�e=���;�'�@�>zROvu{��؎�n:�f���(�Mat��#�W��J!1��.%�4�O ��;)��Sc~����I�K���v�b�pxG`�����U��5q��͜3RiP�s�� 3��a�'E�+�[�9�'sX,��k�}G�ۊ�-�N�Hs���=f^�����"���ER��i�p�>OY�4r�(D�HFjC���nX:�LzYYo��Н�3���y}ݣ��|��{�~���A��}L[t������kP�H�T����/�.&[���Gc��~}F�ື`X^b�T�E��p��~x�W��qJ�=pNC������yj����L�[�Q�5h��Qp��=�%ꉾ�l���P��� S����L̥�<a�SGg1&@7�����>�g���W���z����+�P�7��Ftz%L A�DY�Be{��a��0���s"��{��mZ聿�yu�Y�1j+��������n�Br����ӄ ��wT���n�\�=����6���R�7^�;��k�p��/(`5>7�[��r�O^���䟉��G*��#�F>|[��W/U��Zd[M���U�z�� �
,�n��e���C�(�4³��n�sx�N�8��"{�
�=g�*�7EIf7N_�\c�Mv�5���04��~a��H�YIr�x���h@�\��$�d5�w�/�L�V�Cr�s��@�k�j���v{�ۑyK�:���I�l����^%���*"���uӄ������? Z���C��mj`�dsؤ>
��>�FF�o,J�gw5�� C����l��n���ۡ^ʮ?�F���"�����|�A���R�:�2d(�u�3I��K�(��k����O��;v�ѹW�^�Z�{T�9ax(t���V�
G�/R���X\�Ha �����i��:vY�:Mz��G����zx��ʐ�G̯���R�Ó�E�ݿD���O!M��u��� ����U'� n� �G��N����i�M?�i=����9Um~��Y�c�2��?<Z�o�-4ĥ<���?Im<�������Mᘮ�Qk� ���|�a#��-�C�(����Nޚ
 ��Yt�U'*J"����.^b�*'�b��|�ԓ�v9��Z蚇�O�?0���Y�$X�d�_է*7I���͑���_c
�oWl��k���2XdR<tn��N`���>�EB�-f��)(�,�(�Ax��������äyiA@���d�stGt���\�xy'��!��<hmÊ�a/'k����w�^�91Z�I�I�}w�����H��2�]��*3&����0s���P &�z�&hZE�N�����$r�����A�_w�=����՚T�������2�[�X���9��|�)�=�����R=�#��/�	g� WP1��������ad69Ή�^
%������@�k�2_�%��o��}�_�u6��"�I@���N'q��S�6k��"�U���q-�;���]F�s�7�QYhS*���n����Gr\C�{���X���Lع��mfJ5(e��tJ�4l�2��Ӛ��T"�Ω�2�c�
I���X���-��0n
%��т��8�%��i��jW9ބ��~Uh��A���ꇧ������[3D(�+b>��0��������O,�����c�*i���p�y9��A��xY	�\Q���K�n�YX��F�B�̪�ز��pD�ݴ#As%�ڃ<+�H;�$�2t���
7���[̽H�rƝ�n��ɹiYgyp���(G~D6��(��k��C�UnVJG��q3(TE���`遽�NW�9�(ض�W�W��ߧ�ۖ܃���ލ���Cى�mSA��5;����)L V�����<)�3���k
D�GQ���z�E!>
��4ckfʲ�퓖K5���r�v�5�jk��ns|e�m�R"G}5j޿0��]a�
����`����Ӻ�DaB)���8P�F�Wx� E��]tE?�VpaQ�K}N"�/��-G��,��C9�'ӝg���l��mmS������}�@!� %n�˭6����^�b*�fʴ0c!��4���ܞ��xD;L.�#�`� j^�s�^�*�0�%/1f�6���P�:U���)�r�sxr�9[:C�������%`��?�9`MVQ�	�Y���8W�T�nt��PTj�vMv��eG���� 6�<xDS)�a��e��O��W�?J�`+>Z�D\���F�A����������_�ci�.����:h��2��U�B�⠨�W�i�q��mŝ��[�x�+�^���X��NC��X)���#�� w�c��ܢ��2�	6���ѯ��b�I�����@G����j������5Q$�ٴ���"�Ӥı�;є�d����/i&t�E<�W 4G�(P�ys��Dx~{l/у�
ݶ�ѕg�J'A7�
oNcMr��^Z7*�H�22c�%�=g����k�.���xjW�ꘆ���,�8���1�ǀ�~9���%љ�Q2���]IZ:6s��C ��T��4�$O��A ��O�m؅G�inR� R�vӆ�,Y���w�K1S~�^֟N�������wl�^t���&�>��фQR3"hI�z��J�~���/�)��$��;�V|Vq���4��ؗ�/UFd�i�d���A�_j8�\ٰ��Y_V�����#��3������\�A5��-�72���������£࣌�3?"�\%|(�TWy�s�� 1y�4}ӡ���h�R3�]�y!ƇQ��|���!?DF�kR��)��F��
P��C�e�|�ێu��I"�*)"U���\��.����n���.R}�7��8L�(�Ldk�X��)�$J�^`��k�V6��c�)�gX�E]�&nR�.�{-i��k�hR���;�ք�4����T	W��Q�h{���tX���/�7��r�@S�9�?��x�����#�_񭚤wܷ��R�$z�<�y�&T���!v>��q���(6��JD��),�H���`� й�7��RFnq@ 4M�g������Y>PB5��Ȍ�ɉ��R2,������5��n]ڊy��_�H2^��)���m��A:�-�K�m��]����~��v>n��u��jՌ1�'�!֖_�L/<��=�7�<`�tD���:�4\������	!W�;c|n�ѻo��W���&zG�'B�n�KN}���}m��'X�(�f�A[�y��MW��n΋ph���z���ub����e�܅3w�2z1:#6M�9u^2J5����gJTs�P����Uc��v�T�~�=����PĬ�B��6��<��ް��a��ʅ��M0-�ϕjG��R*���(�\2Q����Ӛ�I>D�RB�n]�����D�黠�L�>���GY>�V� T��2P���Sɨ��س������� �#��m�Y���]-��}z����S��.�˺9 _P��f��nЗf�����Z�~������BvƤ:w�Y���o�F�����S$-��q�9g���$	ӷ��d7�e��o�,��#��+��&c~Ę���iE4���t'fV��r��؟m�<Po����3�g��:��%�8g�VW%���ح�j*������̣ �@mߝ��&��!+^z^�-=)Y���i^`�� ^R3��)u��L[ehZ;c"����9m���޻��@�~8�@���e
�<@��������,���q�d��r��i)��9f���N��s?���m䣌(l��.qB���l��m9kQ���J�����V�i��	N�]�+�_&mA1�׭��VC�Xߌ0nba����>�����A�rw��fW���.�ƶ~�V��2�(
�������j hz�az�'QZu���X�v��}�z��[W-�m,�F��<-{���f�����0e��4&%�*�#b��H���)}F��Cew�رB�N#��*Y��]�m�9,z��я�}��3�uU����w[d��`���=�H:&���2_�GsUw�v6�l�wM���*Gv>��j.x�'h�U)�� ������E������.ݎ������L'��E�v�b1Q����9q��3�i���/ۄHw����i����O�����h�[�!)Am�0�Z�e���H"1�41!��B��C%:Wgl��������X�6��Q��F�>!/._1����_�.�@G����cq���?2�-i�B[j��G����g�or�DDo�wyQ�B��������Ù@�0�t�z�TßU�K��w��ɵ���a�Z�]��Gݸu_�:!�Nu	�t�%R��X�͚�h��ޏ�}8R 9�2Ĭ��^������NN���Y�l��za�e�<CE��z��F^�4Ӄk �y��u�O�C:)��I|��@���� ������.fF��W�����W��]kB�`Ҏ;������l�Έ�SQ�=Ly{K>���P#6Jũ��MPH�g��B��ExNE+_K�U( ��`��b���T��3�e(�#���a��"�O��-aP�1�j.r1m.�lXGX�C�C�\V�ͣ�x��Q��Q�C}����Ջv��v1}��n��C?}�4�~_���_ܹ2@6�=~������	%5RA�N���Ϗ��z�o���B��m���E�@�#��$B�{���#M}�8���|�V)�)�9�׳f�׭<�s�`��c.M��/��	�G.�>��iusmc��G|�_�2��A�
��k镯=j�S\d{̐�����=���\������TxB"�f�����U0�6V���f@��=Zσ��1�Ʃ�!�Ո�8l�!x �]Yޞ�zB���3Kw�`?'�<8����������M��?��x��<c�Q}Va����E�z����o�rIb�*lDA�ٽ(���v�>N%ݐo>�7#Yl�|d�)��m�'�>π#���bn�+��qR��m��~U�&�)^mo��v��]�Ӹc��M��e��ߝN�Q���k��)|T�^�~����5�N����,V[��O� �q�*�U;��&/w��(�tR[o<�4c���,� z��a�)@�ԯZM�f%' 0!$��|�V���Nu����i��^��(��{�ڔ]��jim`\�g(j-KS��$�cz�&�%"�2��Y'~�$*9��`;γ��'�*~+9�8�!��`>h"���ko�	��;�����?L�s]���m͘U��ͺ��C�F�P��@��u�40��m{$�Z�u ���?JyU����M.Ix�~�os�Up��u;�����?��8����=jɘhA[��]�=�	Uɶ�U�ý,�-{5���!6���,���@1#��sS�8��ڇ/�hZgұ�;��i� vL�%3;������Z��|L~L�2Iƪ^�o����bm'θ�DL��Q�x��Q�1{TjX��cT�q���,�щo�s�.ID#ajI\-��l,bٵm8?82d��?%'&����$Ĕ��������++�˳�w�>�ӛ ߒ֌��ۉ-z&�x�ӿjo�?
��0��#R���L�}����y�kI��_x�#OH� Ό�|׳1�;�K��,�S��"���y�ǺP<�*��3��U!������?��+������#����{V�?�ԉEu�1�s�/9uX��QDN(��Y�y��a�'&�C7�'&S`2���*���R���b`�<��0�����4����:�d�����)A�
(9b�_ݟ`V+�����l����.,�_2�MF዆���V�y�t�#~�Y�9��k�G�(<{0%�E�)o;^k���
>nxT�5�SD�0,��jҢ5AZ�|��a����ԣ�T���Q�0���R�m��_�N�E�����@Ѹ�~_2.qܗG*8��WU����y%-'멯�^-�o����MV��Af͠Ê;[�&R���T�nK�f�?��Ա+��ޚ;��Y1Ѭ�c=�8@5�.|�
0����5�D#��Ob�pPE��L<�A��@����y�8���6�ߣ'�6R�=O�GS#�ۺ+�H�!�*f��^uX�yt���V��C%�m�͜ 1�,Gs�	l�
4�eڇ��DV?�e��rJDCۣ�9cQ�b^r�S���`^L(�M���8��}�|���@8�6�,�J���I����ug��.���K��;U�y��o��mp�R�'�D��W{�I��Qy���	3�J٬w��!��J<�&�l����ABiB���)�5�Й�������f0Q��ɓ��n�f�V�k�]2'�݃_����{�'��8;BQ M���ȹ�ﵗ��Ή�v�E.����ڱ��[3)��}��V�)4\�pD?������C;N��@�_)�Ju�t�O��Ȫ�Gvݙ�6�Y5)-��gs��,u��ֺ[�Hx�/W,��%�nEr��T4,}#����+}?�V�,�~�w�˾%X�셎���#�d�Z���!�� �?,�  �~H��8���|�NY�ij������$b�b��ݤ#�[��hތ�wR�r����f�
��J�����W�^W�E�m�}.�صv�P�{.:�H*�0{D���R�cj<�6�=��� ����p_�s��"�x�b(#�2�ݲ\5��\�4��.���L�?$��27�`��O��(�Y����/��!�?�OUFp�����ӡY	��TW2{"��<�S��Zt��_iw<d���W���ՒV�F���khntʆ�r���/δI$�M��U5��SS��s�|؅L��z�ci�M�8��L��1�:�5?j"�A�2C#�9<��ӔL^1��Bj�Ӓ���*�\=��tǁ���t1���q �������r;�5�w�6	Tߊ�?B�܈�68��:g�3�wx�)d�%�����LK�1�*��a�nC�	E+y��������e�-����heo�1���筬	����|&t��PL9�>~߯���u���Te�G��{��"T�ڴ �
�W1�"�t���K��3U�E'����dp�H���e	��W#����#��=J��x���x��4��(�\n��f�-JO+8�X8���d\�_�~�f%`�i���`�u��L�v��n5�	X���zA$�0Yc@݁�n�]��m���uH�m�:�z_2D�
7n�^Y3���<�Ӿ1�9�/�ȭ6�Pmt�1�{�OP�`����[�
�����Ǹ4{�E��.&z>�[��!_ދ�>���dןc������l��0۬BL�z�T�!=v��ҡI�)�#p��v���G��?'�h\�?�jr ��Nc�D�|ʹi��x�TF�G�Gx1���EuXpQၫPJ� =}�p<D��{��z�
f(9G"�+�E�Ȅ{Y&��Y;�@W,��1�s�M����0�I�hGy� ��Z�P�rĢ��p�HdT�����t�Ŧ��,��uf�#�iw�际;j�ޢ9�������0z=�M��K���g�ѨzYE���Z���m��p��}oco�>O{��<��h�R���IX��ȁ۲�X�� ��D�#o�bՐ8�1�����J����^��:��Ż��B�{�z�'�S�iLU�]c� "�;�k滆Ř}�JM
���������G�>����ġⲯP�ڭ:��䋎���@c2R����W��a��̇啷�ld�1�Q��d$��?(�6rͣ>�� �]:� 
���*u��&��!�:�mɅ˼3�h�ƺ��F�"�l �)��w��� 
`uH+Zt'����T�]�����6�>	K����3 ���I�k!��vr�7��,y�Eǉv�(��Q�q?F������I�,��y��m}xiU�Oh����W��֘// �SyFW_�ㆅ]{��7I�&}�:J�����x���{���ӛ��X�t=��9l�ސ�q{�X�G�~��aqg�K�������.'�E�D4��b�Т�R�Q�)lpa	7ȑ�����j�qz}����Pw"�Z�5�Y/��	��T~�����n6dJ�{�K��{c��A� P�óf�J�%�B�w|�h\�	x�KLB&bF��z1<ɇ�|z<��eBp n���PG���A��h|��|w<����'����F���A����P8�G�����=�^�1�o��E�A
Y��E�l�a/�$�;Ѿs��	݌���;N��;�þ�o���g�d������=;���&#U�e��8��l�L�ي��+n� ~ƪ�{H��'4���r��;��2!#��ɏp2��h�$�7�x�����W��#gdu7��������7h@M�(S����=�?�a�ᾫ��z�@p��������`�מ�F��Al[(o��`bǗ�m5kc����rސ)'	׳�*��Bby޼�MEkZ�;�R�<��;O6^a#&Sdb	����]1�*���|m?�0��86�;8�vԖ��s!B�-CR2Hm�F@)�$�9�>�u�^(8Fr.�WD����k�_Y�����AGV��d��?/�30��	C���#�H�iD��S������K��[�kV�t�>�7�3_Jl�T���XF@��p��8Q!��Z�4���sAPu�3��D[�	yojC��-g�B��|@�BojX?�a��[��Ѿ!2�M~iQB���bR��Î ���9|vD�����3��m����}�3�2ϛ�%	��N-Map��� 0�����<j���L��'����$�kmy4I��D��p�w�ղDe�5����=ߑ~�i�|�	��}�f|��9/�<Xt��܍Qn��iO���|�W�t�p��i�6�f�3��!ϡ�kD�e��LD+f+�a1��Z��	{z":˝��7C"�B$X���Ռ+P��9�Lgd��+��'$��oW_�g\� -U�Ǻ���§�B��7&��ʥ�xFx:u��୒�V�6:~F�����K����m�TfŜQ�SY�o�nRdͦ�����L�mg��!��و_Zj?ޕT�W.�\�?�Tgb�E���*}���b�A�2� ����)���d���-�a�0���PyZ:��Ӌ�'ȼ_p��\XϠT%�$]͖5x@�
1K�-vo�ƟE�F��H���tC�M>�t7h�3���q���)�RܹV�`�z|����(ߢ!�A��&�$z�is���}� y :<�G�=��S☋uѪ��	 ļ�I�?�F������&���v�~���xw�mGv�@��  %�U�����CH��2~���M���-^�w>g��;���a�(֑��`��7�D�]� 'r������/Oo��;ꪀY�C�v�d��km	p"��?����	�Pɢ>�1�O�˚�����*(]گ.��i��c@g�`��=]��iMRg?�����4�pum+�cZ� Hڹ#f���
�nSO��e���;��>cPd:=I��b}���^�������E\����$_R��Cjɦi��^��tG�Q��ߒ�3������ ��M֝��Ah�_��gh1�ǩL�����?<�\�5���G//."S�W�UU^vy��㵤 ,lR�5�+U�L�����b?`�f��Y�:.�ra�T�x �<��l���<AFau���`��\������~���O�e3�]%�� ���ѡ���k� z�"P�rA��~ �e�l��Xdl��Fj0�:���>vΗ�_�L���O8m�����}����}�t@�f\љj^^>b���[�MqUE�0��uq�/��.�Qd�K�
�'��)J�������V&V���t������D�1r��Ia_z��E�T��?t�Q��J����S��P�'��"uЎ`�P�%Xi�l�)�0�+���
�8^�ii�lT�����:s��q$]݉�u����v0�BZ��Eg(��J-2��u�
E�{��t%|�l����gn��%:�,�6RԲ~��X{4d/+���
:�[idAC��KyܼUD�!Խ
��kz{��La���k"�s�^���!�K!�(��ߏ������رϿ|�Tp9?0�>�!
����"�I�4�[��XgPe�O����Z̝tm μ�t-���IG�5��;�m����G#p (x��M�VuA���P��3;��a�;��~�A]EsUb��~�>54p�vъg��ֲ�Ϊzn����8"w~B/�o��D[/m*Q���BJM�&�O�]�K;`��l%�4�[O��4�x��C�Ǫ.�3 jaEP����Ϣ�N���@s
�h�Va�0#B?�K��ɳ��k��uk/ן�N9q5��9�t
	δn����Sf��@�3D����E�|I���6�Z���m�F�ƣWh6j�S<�(Tm(�]�U�NS�W�8*�����B�t�=��.��3伦�~e.4 �9�;�ڼ��C����e�c�%���r��J)� v�M֏��kʳ��d��q���@;=�%�N�kꖗ����˞��~g�Si���R��=i��|�@\����.*���])���@�	vux|I��*��D���c�� ٫0���>90J�k�H��t��|)�����JGǒ��m\��L��JĬ+����x�|Dt��[	D�e_)i!V��J�ɷ�-}��ͼ�L����?fq��f`��nm6�o ��Ct(%4M����R�#��3/��63q���l�\���%O8��z�Z+�r�&���ƻ`���; }<�0@�
���=�}��B�v���	����QŌ��,.����I?ް�5}_��)���HQ��&�ځ�%�	��	�d����il:�3�8!�j#����ې�
�0�I;_Zr���S�C�p�kG�k��W���W���*,���H��W����0Z���N �)�ڞ�f �bU���"�����WaA�d�Gu��1�)��|"?ӯB2����_��l��xLfe�Wa��7^G�}G]-� ��%2�'J--���]����+�ۺɖm�������ҧ<�~�P���>�/�k��eS�G�^�*��{O�������N#!���jn��di�@�a���aĕ{��U4���|M���{d��;j(���sx3�0u��M,j|�o�}[��C��M��Һ����9� #�(����N�)�M�Pv�h��l-���^?_��Cϵ1-Z't �4������е�����A�C���#��D�?�n���-̷gy��q�w�j�*9?���<��m��\Oߣ����bM��Ў��<7N�/c��? ��טR�R�B�j��L��@����hB�Gȸ�(L8�����bA���k�`tb�j���^�w�����A��(f�:��d����	<�bR��Z�Vl�t�;�������8�=lx��a��:�SA�G�
v�P������m�eNy�V�&[�j~aL������8�"�:�θ��~�n�rW�!:Ҩ��~d�������B���E��\�r^��fzF����.
 �����!�J����e���N�I�ٔPކ�L9D1*�K�[�~~�ku��V
E �>fd�kr��&����@&��a���J6Nq�a��q��b��.����yE윊�#'���'���<>�W�'������G{����=҅���18�X���2��{���IB�r�)��0yV�ή�y$���~��Q�cc���u�X�u��0W���`#�b��iA�a㺼��M�w���>*8Q�H��l���@���2V��*E�Z%�0�bwH�������%��]2"�v;R�6��@������S,��������k�o�q)dY��k�D��Qw8�V�k�j��V�H��:���6�q\:J$f�*��d�E��D(��|��&0���y@Bl���0牶&�9�mP�Z�e~߹u_[59��g����m�Wm�B_T���i��)���I*�A����.H��I��׳DW@!(�&�/ht��8��} �pl����'<=�rj���;�ǭq.{�5����sy���c�OM0ZT9�Df��:�4�/>\�a�c3;n{Ki���u�՜6R6�_�bW���t�_��}�J}g=�#�<�5
�0�chx���Bx3��C>2�}����ފ�X�x�'|p��:4�8�(o�������K\���i�]B�*��&{\m���x�s�V.�Mȫ��;�y�Z���x���)8�Rk#�vf�yݲow������3NK�N��G��hHx�@��}'C�E<2 ��9"����qjK%I-Q�>[t)�����,��0����������a`c^Cj����3l���e�7�b�"d��>ۨ�����z� o�_�{Țy�/̖Jꀲ�U����j�s�Q����F��^C�ګ.Ϲ�L���K��#�;�e	����i��A[��ǋ�V� |A��ŷ��� �\�1�f��}p2�C�z���u.�T�m7���`3g��6���3g<

��lឰ^32�Pɶ"9X�r%Kw�v�"�!526�(uV��iz!b4�m�Ɵ�������p���#����Jt9�/��ư����Z�B=ct�?jtq��
=�G�^!�ߢ���H��u~�Zg0����/�/|��J�,}юBZ/dV�d�P$��ͥ������X.%}��������>���B��s�^n,�t�=�z19�I�;K�v%����Գ»�@.dd�8��	�
����Rd@�|ۨ�
�#6�Bә���ٯ�,�2|�(�Ч�G�Y\�~讻)�g�|�k���v ��$�h���	��^ǯi��Bz5������?r>��ߗ~�}B�%#�������K��K��-z/�8��ؾ���]���6��݂s;w�/����h`�ݛ
	�j"��y%Ë'��ά�w���G:��Cd	����te|C��P5<�Ɍ�7����%��e �*�ӂ�{#���ݲ@�g��D�m�@�0�3��tI]�\d@U{J=�|"�}@@@b@�Hq�C��u
>�-��B,p[�|=�ɖ`KsN�1L]k_�̼�s�E��;�@'fb�f
1 ��0��KT���R�7�p �F�.�i|w\�.w�S`���j������"g	A|=����/����t\���J'K���Oo�X@Y�Ԓ�<�Ŋ��C�f���2k+�R���+����D����/��KN�t�����c)��w[�����c��*��'�3�Q��{v1�˷jLY��D-�����E�7)ք�b簛7l���^�4�z@Խ�Y��h��.+����P.�"�y^��U^�D
r��ǹ&�Z=����g}�WuNi}�� B�k�`C�+FH�&W̨tbFΞ�^~5K��d���mI���I.�����`yZ��W��Ж�)�&�T,G��9����\�U�{�<&'{㥈e7� �^U�&����ɀ��t�l`��Pڶ���� İ|W�++o�tH�UU%t=X���M����+x��+X�^�;6�}�t�K��0�NC]AV�wS~:�zZ�R��j>�-o�� �kp�f֬�O��#2�~��x8�:L��547�'i��B�n(�1Ώ�M�a7�g���ϻ���
�"�mp�;:!Vp��&O�5'�,�����cOQr�6?���Rs��Ox��w��j��Hk�ma��P�ifi��F���tak��Mdd��+s)��>�����Y��3���"�E�1����^Vyn�*�~�V�H�T�t�Qbx�Fǒ���`����%` ��LޤlӤ�~i�o�]b�d�&�ERŽ�6���Ћ��G�`��o��N5��s*���J=� +(j?��J�v�v��y�F�y��%{˃�EP�]wY�&s|��&���%�G�zz��b}_��A��"��ވ��hb�����h���U�0�G]N�?�9��V7l�qy1�+�6.�k��ξ�us%{� z�+֊�O����o��Fǂ��4��Qd�%HD�h�8݋(�͂���Ή�)��H���W�
cW<�
�$s5�W���Z�t.��<� �� ���t*m�C ��7}�S�� 4~�L��ߥ���fd�k��$J���V��f��1�VIvs�����:x���}�f��]�ۏ�k��q���*�L�ϪH�ݬ�C̞�>���&_�"<Ph���T�Q�����=��~C���)P9��~Q�.WY�JPK����C,��~�T)�;��i��ږ��k�7a��@�Ya�4^Cv���T����itq ^�'pvoXe\��q)h�y>x{3�� ��Z���tv�mH+�j1�f�WpH�9#�S��]ē߾�v'�H��s��S>/�#S>ۊ��Q�]�Œ���%��_�ʹ�~�9{��A�K���n�^�q�H���t�-�)�2��q���Wg��?��1����������ъ��D gq}L���u���1O��V�h�����#�?ګ�P�^�&o��|G�N�!K���q"W=N����+h����7$6��SJ���='b>(��@��84�LD{��w��H% >i:@2�GH���|�11�,��V__�Zh���ȽI;=���*d�Q��):�� �JEx7o�<���b�FG��,�xy	n~�T-�=���\&���69Y���瑈�v��"&�V�5�0�u��e�P7�Ӽd�,���+br�:��ˣ|1|����R�>�f{}��^�e?͟+E̻Ҟ L��*�z#6{>s�u㹤�=<'J5q��s��"ş_[��_�'��&n=A>��/J�lzE��#7����I�F+�d�m�1�]|��C�:֞�
l���?�F"�������2W'�H*I��<�g9@��c�A�=�@�|LWW�Vc��v��J>)��^B�Z07�ȃ�h,�^?{��Z����(*���5�?Z�^$��Q�!�^��6':9YD8� �Љ�D��&|���/�o�)���J�ľ?L�0p1i^�ޡ�R�%�Œ'0�P��^�4��Z9
��}_��ȗ�!�Fi����#.����Q��h��}�!�קn�5g:�,\+�*9.�/��;+4�U��x���
��^��f&F�Z���|�J��궿5L�^Y�5"��pqt�5�0�@�LB�T�D x�M�Λ��J�	��?�����L���a��T��;Hol���H��N�`�|(�Dp�g�T�^)=��'h,��S)
D7|� �S��/��4�Oh�Az��f��1��zs� d;�"���3��Ņy���#9�9VC�-�Zp��O��l���Eu�]�:�-ӑ�Ln�bXB�
V��(�D|!����pz`d�,��LHJ��7ch��L�7<)�*"R�04��P)Ü�^�|r������)>&u8����'�,<��K7+F��]��G|�#6�n8�7����&������Ҋ�/f������� ����f/-߮�=��f>
Y�K��:'r�17R���g��v�5<^-:�Zo�ED��Z��~sj0Ʀʈ2*gӎ���k8ζ|�m�m=7	��c)!�X��w�>��j�1�C�i{�=_��᜔�����4o��2r���o.n�0��_ȳ��R���z�A�m�׎cg��눤��ר�2��>WM�M�S��ְ���a�ɳ;��V�)Q���0���dί%	b�"+t�Tbs9�r��s�4
p��os�87��}J3�֚�j�z*3��':��:�0�y�~��������3���V� (��S(;$�u ^�Y5�>(�i����i
��%��O����UB��q�*��1u�<=нtj����S��}4���c "�Vi���W�ױz�wn�.�3�1���B������W�ko��K��H��M��:�S���ɷpE�8W�"���r[�!�N�:����	D���Y�5�q4�Q5���������-�PLM����4G��҉�t����b��MI'�V5�({�>4��e9t�n�l�j�iZ(���ڔ]�M�0p�.��|m�Õ�$�>e��:ǩ�>�g)��s/�.:ti7��iL�N����-���{�uQA��]�\�׹C��^��b��������.�_.�?H�S�9d�Wr�����F*����	DoM�����C<�j;BA7o^]�y*J��9������f�����`ٞN%�� |Xa�$�F�-h�F�����[ k��$\FI�8��&�s�͖������L�F�VDEX{�R�I�P�<(�Q�vM�@���{a��b��/����NEy�︱��ڸp&�L=tF��1��ߒ;:i��!���!�b�hf	��E�����S!<,g�yDV��>���+`G��[�VUז��T�:��|h:o�鉘
���2sM���-Z��	�������@ВuкN�'��ۉ��/{2Ԕ���q�z{���#l��eiHUM�̧�$pn���A�A�m��_ΐ�ӻ[~|T�;ګ�r�G5Pn�XģL-/L�"Q�ÆK�������G������u�,#a#A��Ϳ������[�����G�L�=�1wm
B9b,4�˹O���7GCN%Ū�p�Y��w���`��̪8^ ���i*���L��,�SQ���a�;�ɯ�$�֜M��Cw�Z��LN�	�.m.������Ǵ�XK�s�"[*�Ќ���}F���˨��)���>��ӛ�3Xc���H�����e�'VX2�%i�]�4 Բ(jQ�Qm�Q龌]{Q�&<!�Ͷ*�~*Jt:m��n�UZ]I���B+T���P�f�a����uq��ts�WB���&O�c�(���%/���jJ�b?�`�d�����|�U��g�ٽ�#�C�w�>�����̀H���Pl�9)�ךY�Z�G�� �����tK��t2����jU#b�S�Vc����4wb�lDw��}��&[a��7���o�foy��v�șK�����A���l!������:������HȲ"{����$��94�	t�eU\�j�YƦߧ_C�%�&����I�����	3���i4��ڤ�Ti�4p�1����b�W|�Q����v��l��$G�?���N���V"��	8��^쑊%M$�>E2o�N8{�񾕦'׋��Zs#�!TDW_g��Ig1��Y�St?Φ@P��,g|�9��)E�ɦ�	s�0كr|���F#����X��̙8�H��W��ߧ\�J�Ks궑/��Y�^���)P��ţ��ף�k��1}vuY��w-l��N�u�،�0���O<0訛Y�}��G8�_�U���ׂ�_�#��}*A�Vd%&���\��E�2^G������f:zX�~�����B��vU,���^&I����A�-�`�I��ֱ0�m	f�N�������/����w���w�`1�y/�*����B5~V�sB�rN�eԓ����^�l��i����S�{�<�/^�sQ�M���1�\pH�ߵ�/�A��k"p��4m='��3ҬL�:��ѝ�9%�����<��4֥�R�pֻ�u��|��/�t8(4V&N�<j�h��B4R+p���ڂ�]��Un5׋`��D��Y���[�̔���y��� �Z���y��-��c�5�E���K�v�Ɏ��[L4fBp�<Q��/o�����+�i�+z�Xv��kjI��ף��-�K���kw~�%���u���b���U�u�W�(�NbY���u�Ѵ����!�TE|�ۛX|���,g�<�:n���/4�J!~��C��bzi�w�J�O������)��iQ��W�x8.ҧٍ'0�/N��x��K�C�a5� ��l�ʄO�u����Qb��_9�u�WŎd�5}������ZO�`���p���_A����2\8��I]�	� V�A�d��#� }�`���rI@��(+a�j�%�t.���M�r'���}I�+��4�&~��=�ӪO�3 $ފ	*e	h�&��F'V4�{��L�3�n��w蔇,�#�l�b?+j��&��ShN��r�ll3*C���ֈ��:���t��AG8{�!��Z����=���zb4�����0C��o�d<=�^r�lE����E�F/{I��$�	�;�X��� �s��6)�x��gʰ�p�!GB�����n�CoH�ܶ���X�Jz��M] ER��r\��X�M��Y�Ik�(�{A��K����Ig�aɄ�N�[H�K�!�E.d�O� �"�����I�/	�$�9���^�;����Fx��z��c���^��O�[��׺i�;P픉�1[ c�9��S�4�a΋��Tnr�J�$ӳ+w����Z�������a��K��m�?���Ls^�����.���e_w(2a
p���53�@����F*M�B����$���͉��z!�� ��G?<:ׅ�k|��s���n�����h��><��r�e����!w#i,���t8ү�r���CS�e� ����ɀ3/h��-��0����0	$
�������.�C�Z�ֹ٩Y!����!p��'3�����w3��D|F��AI-�M�cx��Hʝi;���g~i���R��\��t�z-Rw�����/�Mܴ)�$��̓Gfa%�ك�&��h�x�n��zc����k� 0��QP��	Ra��I)�r������l��D��v�{����@R�L����^�hˆ�܍���}�cTH9Ϡ5	*0�-���q���"�#�A���R��\z��>�V<;� �H�ݑ.8)����núZ�;�M��lY�Y�ݨR?0�
˪��1���=^u��}j��eM�+<����j��s�v�7'F�:q%���&��LI�j���v�){��#����內(��
yY/�S(�L��̋G��ci�T�k�S������\���G,�YO薆JÀψ)�aH��ob�߭�+-g���6����g���L�A������_�j6��
�&����bf�c�j� -oW�e��~�A����p^����,�~?W���?�xR����y�L�r�.pi�lA=v�Ģf�RBQVa ]_���E8�6A�Ԅ��%>s���}��� ;����'�ߏ���T�w+�F�e�C�ӕF��1Ћw�C��͉��=�$������_�+lT�=L)wg�k8��*�Do@�Y׿��OP�l뭱5�Gbϝ-ƙc�����8ܺ�N!O�_u���]e���6���l���@#�kx����]�g���
6�R���9&<�^�B�� #�Q�Q/�d���S���!�s���"�}Ċ�ɔV"�\��U�<�#����?8�Z��5��l�&q]�CA�n��y�g\�D#��L6�)I�Jk��SBU*�3�_�I����-���[�}f��Ҧv���J'06��Q��A23i�1��-m�x��Z����:2@���\?�ʗN5��`����iڈwM?��"�+5�zõ���q���_�3�pPvS
=h+�%3*W��S�tm�+?�O�br�uc*>M�j�v�i��Xٮk^[&�h��J�Π�z��F�)"�΁)����5 $E���|��P�͐���������_��1ӳ�k���̮���f�=Ǳ�X�EiQ�Cɦ�.�Mȋ7�o�v��R=3鴨設�^y��J-}���T�lO�tˇ��Ɋ������Y��<5,^�%�|{�8�|�&�7��mFz�G�9%��k�h�j/@2��F��W��I�j]b)���ߓ
��7EM᧣���}�+f����T7C7l-Ü�rWNL�@�xo��
I4^H\���KD=���ֻ�D���ز�g�o��@�փ(��B�@�pXb��-�z���g�_�s�:�Lϰ�B�e���V[j���U�EA�)�
��txls���P(��B�x��fA�q-�M�kҩ�rI���8����
s)�T�E�L
�FƬ�q�x�t#���Q/$��<��Y�ʍ<�*��cDCض��rj�D�q�tn)+�����	���V����<~��5���L��H���>�=��'���|��o9���v�*�3����/��u��!>:h����?�X���+E�Qv�����Ʈ�T60�'���֜:3lv���2ؽ}����y�C�&�����Gǁy�*��VM&5t	�Iy��d)���L�:!���m�i k��Y}2`93�kM��:H��{�b�`��%�|��@gk�"c}zq�3\~-$ltP3� K+r��bp�2���.�l�a��+޶ �<m���X�Zy!'�k��䱲�7�fAr���u�'���F�N-hS�Կ.���L�s���m{'���Qm���D�U�&��������&�x@��c���0�(������aT��}�$�$�f�5+�r��/喹��Q{��m�W8��KF�����o[�ԓVxs/�"��������K�YZ5۾@�(�n(�����va���-&���)F8ßI��+��㶩y�t�s��b����9��G����غ�ƪ@|D^jiD�ң�I���,�ϭ��kx�d��OM����������� M�c��	�ͥN)4>Yp@��P�wB��&�P	R ��H-��k*N�<n�@Pb���?�nLM�3�����*[�M�'�/ؑ/���[G@u�;s<������d�
�������m`��5A�P	�kI��o���!��X�^f6�J�$�K��.����2)4x��uOhg��-"��9xN�+\M������vY$�(�Q?/n����4�����LYBtb�v�&�ҁ����&�t���!�K�|J�U���Dp/��	�c�����X;"�`�<`���7aL"ϝE�6���7U�&���a������E��T#�^#j��M��ʇE��?��`mM���-�V�\O9����P�~P U�ވ��})(��R�UW���ZG�Lߤ��C�X� x�kb�^�{��
�ak�l#eM�\�^�K�ol o1�)n�����I��k��k���
Z�M?B���#��I��I�8�b[�@�,����uM�v�{�g��I�H7�xϞ����߆�v�S��J�}�j��O��b�9w���W���^�����9lT[V���]� 8Í�3���Z��>�%�,�ld�˹0��]���/�����|�-+?KQ�l�0AH�$众-����3Ȕ�ל�����,����:�x ���\�-�B"[B���Eh�l~�\@윍e�j�R
=vN�Ms�D;��u;�NS�3����љj�E��vdߌ |�m��5�D��f�/�)=��\`@܀����Q�?�D��ѾM�G�(��n��� \�;O�^ 3m����ED�?��P�;���Y|4�k�u|���A��\�N���w/n|
�%��ާ�kj��Y ~���t��Ae�I�2m:t�\s2q�Lj����5:�Tc�@�HoR�\���V~�v)9A��=L��^)e1������{��ݡ��ű�۷t�è2)�¹pEbo'��y#Vr�c����/5Q<�1V���au{�>��O���9`d�HT%��\���K�Zo%��9��y�$�8l��_JPR�XJoՎ<����2���1'T�ȡ%�4�&���Q.�H��qϝ�� �)����HU ��]%�9��<�3��CD�ԤY��O�Ӯ�1��J(�E� EI��l��Q��납���ٚ�C�P��P�I���q�8��l����x���SV@����[�R��;ʬ�۝^! ��]r������:�D9ɸ�2�\�e���܆!Mu.��O�we\�G���t���Mlڌ�����F�]�N� X*�Z�K�C�s
@ ]���#���@Y<J>{�)�@�iwdW�n}��E�zt��\�5}�]ij��vO��-hz������"��c�p@��`��A����%ŧ���с߶[���#J|dmC6;H�/�pTY����þ�m��f2nS�����+�b��n��@��{�kn�76��N��њ*��۰��DiU)�5k�5}f�̨�Prމ�;-R?�PD�*e�0����:%^�3U�.�N *�n���s����))o�\�YtF��g�h�h�ܻb"������R&>m4���z<����v���m�	���x�F�5C9'Y�A�L������%]����G4�	��]��1��驄ǗJ�g?��ȜZzd��'��X։=��8�n&��q��3Od�����T��:�l�ͭ0!�e��@�
4����m�z=��˕�	kɋ�ʓVK�{O��2��J�@�<^�>(x�)�ώ��лP�x��Y�ļ�wN���0��.`#��$,tU�(��p����S�"t�*h���`��y�+�\p�p���m��)X��y����sAN
u�(n���[������BB�D�sIF�\� `�`;?��s��������S��!'8�ˤ����)T]��j�V�?/��&��/��Q���_5/�#����>n������':��Q��M��-�Cޯ9
ɟ�����~R�=0E��q��ܺȧi��i�5Ԟ�:d��,Z�ˤ�*�г~����|M� e)@�1���H�@>���틖P	�t�M��q���
���hTD��V�Q�7�3()��,�)A�h�̶s��5��-x��&bmz�ڵoSc1���g72@�����F1h���>��N�<%�4�~�Bw*����2wR{2�u�t�k�a�<�>���T��N��K�f���T�a�Y�O��Y�^��ZOh#�H@O}B ��d?�D��U�iǖ:	ѹR_�1�,�V�et)�!t@�8���<�" 1'q����0Z*�����.W�t�Q}
�+�e�G%Oo<�4�=�u<���68w��NbG�o�H�9J ���fHiu���ʹ ��1�a�g.#�w��i���M�� �+,��2���j��\[��H���x�HԊ���8���ׇ(���������
p��Wu��z*�:��%f"�
���;�mryUni����@�q��'~KZ�@��P�V�u��(�Ȥ�E�~�p�}�J��C0,��cVVk4�K��*�1���q�-�v	W}��>�K��z���� �!`}�o��Pe^Ц)�ݦ��n���Fĝ��׍�蒶�-��6�YI/��>��HaKR�s�b^Eы�h���xC܅���&ˎQz	zI%I��L�Z��S��<�<�f��]�y/�(\���!��+c����+�ˠ�]���n�|��xx��o����9�8H�0t��o�Q�C�7qHE�%t�)I�PvC��X�S?��@M�-���	�я+a4�;k���@����-ol��¶ g��>mhZ2.�â��I	��ǃ~ɒ�=�������i��_tq�	z��#�+�z�:�u.q�p�n)�<��!?!��?�*`�˸gY�_�XԺH�epc�e/�2t�V��%X1$��C������ y Hs�	V��5P�_��Ӗ���+%�b;������5���T\�B/c�ї��
'}&ě���i�UZ��V�#ȯ�-�`QGO�C����-.��X%͔9gۭ��B�#�]��o�{_�oxgK� [�ʀ�"� ��n7CT6k���9|}��P�����p�W[��7[�X��i�wQ칀���َ�'�>�}\��pOf��z+�GA��/�'�\`5�e���e[z;Ǝ� ����x�G��N?��C�Z��פּ�d׎8,u�=G�ǐDh���o��;�8{X�g_>������e�~�9�Q��x�Ȼ��;nW�t��թ%��t�3�x��8՞�S��ܧ���}�	��=�u�2��_���G�K Xɰ������E�U5N��}��z������j/�20��䐇�B�gQ�,�j%�&���V��c*G�/!�xvjnK m����x�)�O����z�z�.�Q͏�[S	���&�{b�O�Xqh���Y��} ��|,�$�.��Ũv����O($� �p��\z��FZM�lՖ\Y1���T�صラfâeԊ��kZţ+,7��o����>���Nڨ`P��t��������΄y�@���&��������w�D��r�aE�q��r���*�Ӧ*�,��X՟ߔA��r���kĒ���}�?9N����Ce�¾����W}zma쒧����i���|e�{3����%�b��z�)�%9(�s�0z���@eO�	Y��垑�,p�?*�����]�˒?�l|�l���+�6�}��l��ܐ��NF�gBQ����5v8'���b������K�ض!3Y2Ikg�y���|�bk��G/P��z���G�����!��N;�eei�E	�BJd̺�QT�n� �]AK��}�qe�Q=vbwj�7D�#����;��RI��f� 0��v	qokdτ�$���f��!��6��7���z8�����o;�X3�NRx��ի��*�B26�<'��:z{> Wh�P&�W=���}xQ
1#sCn��Kf�A�E§��.���
u��FQ��c�M�������n��(4�oa��Y��X��4K��0�_�On����XY�oO��m;9�>M�[@F�|����[�`^ ��+l�d^�Vڤ�U�c��L���	pC~�mԆX��T6��G��/�zAKĎ"WnWXdGTl�u��tgK�-��F��)���
�$�ԒV3W�)��#���5�Q�#y.��a#a��/9Ϥ���.�_lnb�-Ֆ���҉�!-�I}t�+K�6a@$����)ff�!����ҳg�Fxu�u���O�{h���j�Y�ȋs:�h&�L�{�(	T?$��~d83(�6smൂ�3T����y8U,:c-V��Wp%d�(U��Pal$��,7D� \	�c���v�j��ӜNm`�/���$W䴳"���A�$`y��,��@sy���5msK�FV/��s�K�HԞ���2��H·�g���_\�g�"�v�]ǯ�����kC�a��\��CYn��B�f����FH�����3efM��82Mϟ�[XƢ��OG;S�c���h�^89[Jk��Ǒ��"��
�4���^R�>3Vo�%M#��2.��W�u���jjvZ�|��
V�k�O]P�EQ5f����{_gc� $s����"�����<�7���|5�Gaف�����
��{-��o�����>�����.�\�I?�@��0�U�_wlR�X��P1Ν�f���^�a����X-m�[s�B����G��A!�� ����r�@�?�u"���w���.L�(�T-k���0�(���%gsR'����~���)_JZ�^!�GL����p@%dX:�(ш�R5Uk�ysŉ.�;/���5��Bq2��m>��r�`�o��IQ��f�1��}�ĕ@���Ҙ���֪q����募�����D�������{:�][�m�Yr�:������ 5���Ѕ�T�(�� `g�<�'�*@@H�7���k��И�@�ǯ�}qL4�p�_,e�R�������K�������|�t����.��N��Uc��e��ޡ�m�@Q�0N����YZ��6a� }ʛ������Z�"Uƹ�5avܞڣ���+����W�s���D�X��P�ؑm�p@�e���f��N�{��.���f>]$F(�H9o��ȶV"\�6X�5����8�?
hN����h����{us4�B^��r֤�o*�P}drr�G�b�F�z��u_�G�0�l�G�4���c�vY�=!�i�cK��3 �x�!�1�[f��Wn�������'(z���;��GV���ZǟN�}ӵ=j���A���='�)�`�6��Lg'��'�X�g�$O�Ď��}�Y:�{��ǩ^��?@�0؈-g��m�d��)e�^�����c�-��y���%˝��Hex�=�DU�|����M�Iͽ�&�])db)�Ud�Ȁ0%�v���UL��5=�I['�Ճ��^1m���ћ�+W��GI��6J�HTc����������S��	�T���q�*��P�\��P�����yO��X@P�GT�-Z=>X��p��X�ɲ�Dn<�����������5�Y��mE�_����kb��Ev+�iRI��Ns��i?6̋u�g��;�dB��m/���x�Qa.iw1�����o��FȚ*�4ݫ�`;�钣e-��О��xv�jᦫg� �>��[�����CD�s||)���ށ+-ʪ�Ab��4%��0G��"U�������Gg^$�*?�ذ�t�R9sa��H t��8����@�t�4	����������|%�;�Շ�A�w�V����C����#��'��%����9V ���,��0��	S�_u#�n���]�sMoW�(��Fr�{�Z�f��!'�c]�0��UIuܥfK2
��+����w'F��hDߙ|�WP��J�e�_�b��<���ؠl@ <ۈ�
�Lv]��fbI�59巋�}?��2��I�j3G��x�v��Z֐�&� ��G!t+�hU��7�LrZ4֓wSX� �;���
�N�/��ϦO�0�l�g��4�n1ōN���Ʈ�1���k��&����Xv�X��ocO��!=-?�S�B(�oS4�4<R2�������?�GR�l i~�C9%������N���4k��SDխY�bE�>7�������}�x���j�GBf���J�G�"�{������r�+�pUܸV� �ˣ��*��*�C��!���qa"5��~<�&�&Sz��Z��[!���_�sd��~�C�ҙ��҆�h�)qC�T�޲������݉w��a'YV�=��b�	�6Ygs)�A�Ԥ��m}83�+���l��?�݅'[���GP����B%�	��7�;�ڥǮ�a��_��.����cI����U��3.9B\�x=p�7�S�;��gS�8���b������9�XY7�L��P��JZ�����XE��}l[���y�PoO�a� iY����N��@Q��0 h��_wD?�V�T�������s�I�s�+��C֢Mj�mw�I	=�Oů& A[$��Ց�1,*��a�/�� �3�^���ܲZ*�-*���b�g�[@%�]G3�e����v+��lf��l*���o��Amf�6d	N<)_<�`�u䶍�.�V��R�T�>8�oHz*G����z�� �j��}�GM��{��3Y��ZlM�Uaj3ۮ��mT�۩���Ϗl��"9"𐀩/.!��`4����}~��#Ai��ÄҪ�<�w&��&��aU_��a����D�[��g��΂V�;i�����;��� �!hnKOF��֫��7L�a�\����[YF:�v+(�rt����W�S�U�Y��-ΓT 6����v�@�KtS3Ul��x��w��s6�4΅SX�l0Q\���@���_�3M����i�e�
1���N�Q�R�1Aѓ`',�ɈP����m҇tWQ�)2�4!C��B�~/Y��/0��^q���(�̣�Be�-bڧ�r�]��/�����ۼ#5u�R�[D\k���MHN��	���9���4@�46j�b������b֍��Y6V:���`߼֑�M���'�1U�Y����3�V\w�Ǫ�l�s�V� H�M���V�B@?H�_нb��F���i��FEg���i�{џK����
�5H�ꘊ!�muyF}��Nد�f@���aQ�wu�#�̡���^�L�"��aX�t;m0x6�	|+"M3Qs~&c���u]��R��k�j`vg��_XtD�)SS���eg�"��ʏ��ƴf���vyɳ���yc�6���\p�@Ky����@�~�鲺($̧���(�h�:�Pp)s��0\���i#nY����v[ٝM���O��Z(S���ˍ��uL��z�f�؆���y�ë��pu_��� �*�jH**�,�����ǔD6}�lRI�"��k5q�Ms1� �=n��+T���N�j�����|�`C�Vuv���%;�(�1�����nU��1Gz}kD]��W	F�F)��ћ[��/�F~\|Р�
%�]j7.x�k'"[�
N,��L~64L�=�IO�y���&�_��;f9Z/���6_���E]�O��0;�)�|�$�DF Ɗ� ���`��#BD�R��_�ؙ���Ԧd��[k���$����� !�Rwe�\�y?��pOe�ǕR�,�M���ef[�a��C�>��ʊ}<�bݬ��l%N1�|��S�W����YѰ3�G��A���fb9��dC)a_(1X����H(z��#��0U���:֥9��ť���<M�=�Z��:*�]��}rd\���&|.C��mUw��x��DJ�B"�F�k��yu�G�EJ9r����z�D�x!r7ٴRO|�Q6���M�C�J���X��A,О�Y�1\7���j����=���j����k2��9�֏j�����(��/����g~���L��!�J�[���=ƨ
������n��M{�8HԻ�f�T|�@��
��(.9��̂���kd��m����і�]���MH��Jn�MH���9�,b&�*J��E줁%I�ɃK;O ����l�YQp���}��_M�� ��o{�k�T� ����hl\��~MZB�zrn���p�A�P�Xh��JD�Pc�?���ְ��c P]?]S�x:5l��M2uC<�hI��eP$�<2�R$��ٚ_����c9�m �C�O�k�t�j�
4���2]���Anq\���8��ьsZ�Bl�+���.b�&_n��B;L3�γ��)N��+}��jH!V��c��a#{	xk����w{us�_�b�in�ٴC�~�Kh�z�!��A�-��B2�"p�9Sb��eC�瘧����LO����6���O}|����1��雎j����u���lƷ(�d7��Q��^�"p�8'�1�" �)u@<��Ԅ��`Y39�=^�#�v��=������J����E>�kF2���τ��X�@LXg�!�W��9���҅�ˍ�o��ŧCc�\�`)Z1{�uaϒ��V���%���w�C%��AIiˎ/��:���Z���x�{���[v�g6W��\���YJm#,̮� �����T��ǯ�O"�+�����Q���3�sk�����H���X������P�Z�q/��rBN�?\ߣ��ԥkQ��iu�E�^@�o>��������,�XGpux����,:kpߤ�k��_
�����m+O��r?�o�A��V:K*!D �¹�{���8��o�������9���vA��w:Hd�%,�u0�®�F҆S9:��=��?^ƽ���ӽ�V+Q6�5�-�yؑr~�����i��a[�on��{}dm���<���s; �$�G�,��==�9Fl�3^3#Sp��5+��{��������Zn<̡{g
΂:��ގ���viec�ыk��G�}�rQ����Psg����^�;O9��^/�[�56�N�^ό���Zh��B�s�Ala,/��I��\�����"�u�ϭ@�Z�M�sӜɐ�����0�0��C�����5�Pd_	e1/��]�%BP��"��@������@{��	���V̛R�\>�w?�N���5�+m~��M�)���~�{�r �ŉk@^�Rn��4�dڶ�>aDf���F�I��n�.�P��t�d��U]��G����X;+(�;l;R�Hi�V��Y��cXz �#���d�\ǰv��B�����8��St�r��h�m3�U�O�0^�R��(b�U��^ơ�3r��0�Mq��/�Y�U6z\�!O$2ʝ������u{WiP�Iq'���: ՚����A�v��d#fKD�̋	_��b�4yw��M���`�2�^3�`��TfH��	�,�E%�;̲RȎ�R�(�ؗ�eq�%Jy���÷7��I�g����:�֞[07��kk"O��q��t��뎂�m�u8��M����K�&�R ~9�M ��_���}��Ν�<\Vא7��͟���B���Z{�/�^5���d�L��u��Z�[��F�
�� �M�&�#�P��dۥL[) +6��c)?���,N͓{�x��j&�A������i�0�M�C�RKa6��Z�a����-����>�l��+��	��cM9c3�9�o�/��VfZIx1��m,sw}u��2ݖ�;��aSP��z�6@~��"X�gߙTL]w��S�Ss�+��l�GG0����,�g^A�<:!�N��?7"��FS	!B�Hp�=DhQ�n)��.̭��D6��<��3n��x$����,���bL�y$/w�*ڰ�e�ϑ9�C�`~���sTI٣�-�T�"lc��13v��!���?�[� ׽gH�p*�F�Ұj�D`�����56��`��X�	�ݰ��q':�x��pi��&��1~lW�__Z���E� �8�p\���
�uBu ���oPP����������M���Kؽ����:8naHz"ko��=Fӵ|4�CJͳ�p���R�VO\��@�s�=r� ����q���і���گ߉���|k�N�T! lE��N/Rp�4�Q��ǡ�*�5��3�N�2t��/���\߰5h�/�j� G僌�$�ժ�� ���PU���@����o����kA�U*C}ɠ����!��u�5@�XB�|�VDl7�[@,� �G*}�o*;&�˽���ȡB�h��ʚ�{5���g��/v�����%I7��{��!N)����&�㭸A��wI*6j�6g3�I%���c�����xYog'P����Ԙ6g��m�U��5k��(|^���} +������:E����6ێ���� �lN�Լ���t�	)�֐`��<�� �M�H?���.�˒�`�3 �'�l�x�n &ss���$��%?�>O���J+Kh�!�|���Ѱ�t�,�o������a�u+���`�� ��Xz�c?�^��
zL�IL�����3
yt&�+�������?@ yY��hDD.R���'�ǧ�ܐ���+`ǈB���>��>e�b �T�ڱ���c^^�u���ݓ��)r`@=Wk	�ih�8C��JY�N�\N�&�O��흱��f�}g1�65�A`��RwaO�Yۜ������?��K���+���7��(md�]M�0�O�+��ʂ)	�7؁�� �6��R}SV���.�y?'����� w@�^59�F�
�.�`��;��y���_b�#f����ȥ��PD����w��`E�����p�ȶ���8h��j���z�E7;Ҷ��0;�1Y�'J2H�ڴ�^<��u ���	���i|6��.�sf�n}0�`�|k�!L� ����g�h�q�`����\S�'�������2�, ��N�ʌ�q ����Df*\j���~1�a�}��ǘk,���;V������Pl�}�xwb^��� �Yϑ�\���F'�(��0e�Y� �G tm��w�2��OZ�����,����5H�HE��eA�($ئ�?�5�~6)"���t����FrnrA����T���P�l�J�����-����[>�L9�8�+c�q�$�;�A���z��������R�QiܘzIe�D�M񵐣!g����6W�Ejv{�Jb�	�P[����-��b����o�1>]>Ү�)�^��;<xM7���;�}�"xP�����6���"	Wۢ�ME�{,<S�����k��D�HV�(�b#?Zm��� ���=�̖�^L�"�� ޢ�` �*F��Y%�&D[LL�������~���u�(�F�1`dN�e,��r���8 2E�I枞�c�7�~��Ua���V3A�n�~��y�|Lb���۫�4�>c�c(v)%0�{�ܨ�-*�9���~'��g@[Py:�}��ݣ�&��*���f8\�։�0bar�Щ�P<j]���>v�q���W�bcq|�*�j�j`�"�sC�;�huӼ��p0>��j��^�G��dZ�h�G/���B�m)�o�US惭J������4y@!~UG"��'�K���a5�ّJ�%�k�y����R�W�E�#Y$aR��XLns^��
XWHԒ�-y"�n4�X���b���1��h�B���4�]$��1��5w6,��#0�@X�At� ł9,�m0��T[,'�|����%wq��L5�(R�o�ڱ���@��zU�q���BZ��_��
�ߘ�VY��nj��C����:'��{�>IFXB�L���&������A:,�‽�~�����fVEm����qMІ{)G�%�n�#'���|]F�#w��I�K�N�1L��8���G9n�NW�+�R��_��NJ�:>G��@� �g���=�v�����&u��\�����N�nuY/�S"��Sp��U(ڷp��.ʖ�y}��.Sxf����O���v��!ylq���ID��I�E��#����Q4��40z�^��-����r�
�ʰJ�Sa7SD.�i����Xl.�r��{)�*(׼O�ypY�M�-��X�BE4���r椄�c���@ϥ��n5욚�9�E�w=�B��H߰Y6_�
x��'�����������DĹm �Y�=���.���X���'�,���@��q�j�Yx��[��ؓ���nWj��
�y������̮F�&']�~�����#�Bn6*_��^:ǖO�4䄥!=E\��8���w[��`�W��5|G�M��x��������r�k��u6d�;?(������ݼ[�V�}�Gx�13�f��N#���8���@����z7->A6ϵ�� F���3jh��z%o�����.���w���\%��̾Z%HY^�m"�m�a#��]��1�YŲE���-���?��g��T\��:I�Xn#u䣢�k�yIx@����ñ͍e�"��N_nJ�$m@�B^����4� =2����&�ݼ���-ҝ
�ܐ~&�aĀe��s8r�=\~?�j�e	P�$dwE�e+��8![\|�q��4��TV;B��1"~�w���Vl�7��	;�1}!BD%\�o���s��c*�)^�'�U���\���K��.UC����G�.�CW�':e�'nO�dg.ݳ���V��yK���E\3Y�.gpPm{RѝG���y�-$Z��c�X��8�X�⚑��U[�&�5�I}�)����/��H��O�+��A���g�Z�`M܈\����|��<:B0���B��9���Zx�R��&��%����F��]≢@�{kb_��U���w�EE�d�eP��xn�9/s[X�I�Ȭ' fZϲ	8�E���=��my��~X?&�!�~=�e�"=4��L�Y��:��sQ����t�>�J2��C�&�����X����Y�}�X0_�+��'�%f�=�(�896ò[����s@]fT!��B�ǵT�m$� JԔ&CE���K�N�z���\x�MԀ�Q��7��
%�ك�L�%�a����@����b�r���#S�.��e�2��"�8�_�v��ge��ѠG�͞H8�%UT,i���p$'�G��5�w̄�M����2T��'�9�.]` /��Dg��J��_���7lp�����ܸ*"��s���;'���VrF�jc�P�i2����ub#�d����
�m���NS��]n����[��>,�O�I	�L�D��l�u�D/�@l�g�j5���Iڝ�B<��_��ʘ}~J��jbFp�Ke���60Q?|�`2�S�C>g���l���Ճ�C.q��R@�s�	Bt����s37��_�o�;�kH6Nߡv#������-�D�&i�aZ'eZ@�c��$����U���At��)kE�*���6�Y��K{Ge%	���>��*5C���a!�z�5u6��(��]}v�>m����߈�;�f�yυ;[Ɲ��mt�C!��|.�*:�zZ^�6�v>"q��F�R3F�"�5��	��1�0���!�[b�'S�73/#���Iѡ�oN�U�?�i1�Z��C���$�����c�֋��b����d�q�Ɔ7��XS�&D<M���ߧ��������л1[��g�ԴƋa �ou����+H�:�tRʏ0���VSXM�$ܨKD�2�P�Ӫ�a�	^.��,C�L$�t�l�!n��!��O���m�Ҹ���h�Z9���a�w�ws,=d)�߰4z�ЉQ:T�1/o��Sp�4�&�+�Uy<B�N�;D����|�jW,����av��P������r����B���0�mn�>=>��h)���N:����m��]:5�9��|�?�㪩���X��< ��cW���Y�CR���S�H���z�&��;u���x��2 ������_�p��'O�9]�.�����Ԃ�Mr������P�y��ؖRg��N� L26Y߈DIJt��uOL۹�a�.=Ź�m���cs��νf�f�O<5'�_ɞJ���W�͂[�u��B��*"t��g6Ȭ߄�7�6�f9mM
�d��}��Wg�+���>&z}0��� 0��h���C�ƯG�i�"��{Kj<��4!s��A��������.8�PwZsH:���,�kV 3���t��+�5t'������3���$�8����.LgZ�u��/�{���d��A_U:jz��N\���K��La��JˣX����h�o�/��߀�fТ|�-`#��'���o��*��ڒ��)�޾�F0��HT�X�e=���Y�nY?B�Y�=�ۙx�>�duKy)X\�U}%n���WTE3��ь�[)��+�^i� �X|��Ƹ盎2؄p���fb�z]����r�Y?NB���9 ��-��Y�S�����åM�&|�=ּ�r+�o|����UAs����;������VQYP�������ex�vQC��*�W*f��/p�P+V+���٪�\B���<�JC|�k7�k�aB~K��;�`щyґ����/{->a|��5��S��nEf����.�ǜ@"�О'�R�񢠃�f�L��3߹`��I��ot�"c��U}��B���	|�uظZe;�e	@�z�ׁ�� ���n�܅��h���L�>l�+7��M )�Bc�ͧs��un��^����]L6�;l�&���l��͟�3�2����a�o�[#rjbH�w�Y�l@����=L����m�����J������d,�������|*wN>���9h�TG7��24����[��:�7�Et�g��vs�M ����7��������Lz6�=����n�a{& ������C*M^����5Pc�ݿ�L��:��'��2�����1�=R�4�q,��k���7���w`h�����l�TTq��B�k^e����@����z�Mɰh������:����Yp��i*�C�]C��V�-�e��(n~�b �t��۲��:(��1-����>�Qb��R`|�5ʙ����SmR�D�g$}O��;�g�24�M~�7&�s`���h%�}ʬ4�H��2$)���i�C�b��ȶ���l)�������<�`��b8���r�UU��ձ\��1S��T�'�Q0�2C�� ў� ���W-qB���>G�Tc'������Z�s�����R6N���|#́��ubW����s��~�6;���py:�*>̹�F?Og�Y=W��
腂~O�ۼ��_�@5��yIbo5�m/T}�֩j�*���@�>��+�s��X��,��8KڀW�:�+Ȟو�~�I���^���Z&�H�:��]ѹ�22/"	Z�����>R�@C����U��T�D/>���c�@����o'�5��a=MK�Fh��?��l��F.XV*���V���h�	H�:�e	:J��vT�m ��gm���|���>A\|qRaK ��(Ω����>�o+�+ʩ1@aLL�U^�e�]@�{�I]��!l�XO�,zc�}���s	پ�&�
����#)J��4�ԙ2ȥT�@C��v���[�j�9m�>A~ɐ��4��m�L&p|�a�Ɲ��޻z�ymI�9����GCۀ1ռ�����Y���B��/��&����A��f����>�;�N�i�q��ڵ�'���uHr�e�0Y�3��`b��fK�R3�s^Kv=�� �	��ƍ����e�+u����-�^�F4qM`w�2�;*����6_^�M�N���_�f�4c"��|�esvL,�-����r������-�*�&�s�Wy�I���i�z� �v
!�!E��[{\��I2�F�����n�b�)E<�͌�:�u���+��fV'�I�d�&��i�f6��Y���Y��~L2���4�=�]뻣�1��$s�Z�B8R#|WLsX�kYM�_�C�bZ�~)��ĭ�]ʸ`I�dI#�:fH��pv����<� 4j�����⡏/cvH�U#:x�CYt��B	n��p޶��x�M⩜�ȼ���)tlr���q�ץc�۲��T�Kw)�r�4ۖ�fjJf����̘I^��"踄���v=4C�X�:�nE���;kx�"��w��a+�H~Wܵ�'��ǘ�a[u �Tk\ɕ���p���������}Z��DFF؉ם�r�� �"�����3�1S���2z�W���OIx��c����K��PD�~�}&l��0N�N�A�ӂ�g���5���T��8�����ާ	����������9�$s���^ԣ�W�wZ�awp�Hw*�,��j���[��zqM�n'0��rRY2B3���D^^	��ڇ��.��������駜&��q����i�%s�q��߱�bz��xȩM�7���tT:k���}��r�+q�6��wZ�"��tt�E���6K�ࠧs�ш7Kp�=�vi��ܧ��2���AF�X�hG���%)�XqVa6��M<db�~�.��z���6�@s�-�	��0u�C���$��$�f�635@s!j\���|����I��xcQ�d����Z����Ǉ���Ye���`��*=�=z �iYK�� ����g=*Q.� �^=L0��&��
uN휴���| �r�#T�W.�^mΪKD5�)��N�MG�RPC�~�B��ۋv �-�����X�M�Y���*2%��Dǔs�
8p�{L��=g��'�b=�G껇{�	�S݄$��`)�]���Sy���		�dƎ��'U�͕d�5�C���'&��1����G��Z-_[��#{$�/�9O�����h�����h��\�W�%�����/�$HemJ��#-3�o��rƇI�[����N�g�shg�<.�ra:l��9ž��r3�&a�J��k��-Y
��)��2���a��>�ZK5��y�Ć^S�c��~����7��b����l�B��2��me��Ϝ��ƕ�HB9��WL��]VG�!�����#L,f�s�B��@uU�w29N�-(�*ݮbVJ��\O����o޴�|�_S����C����7�&&�'uצbD������]����^��_�N����F�N�?f�.FT�|{⋳'n��6M�Ҍ�#��"���8��l����.�V�N���0��_��MKy�ğ���f�>G�t��ͼ>�5����$%�2�jns%q�V��Rp�|�IR�]b����r��/G~w�eέZ�k����|WR`���o���.����0ޏ/�})X�@�������]�!��ynz�pY�_ ����IU3Q@��ȯ(�Z�X�gW��	m"�$hT�`u�\�,�����\&�#��&Cr�N:�] ��u�z��A$�N4٠��Ĺ�,� |.�v�GS�ȴ���l6YE�<{V\�2�F5ksŻة��%�n|H㫏��fA��Ѥ��J���,�sl ���){�E��(_u���x��0��b=�2�z��d��{�|��>؀���(���Uǖ^���=^���+��-g���旋�>�1��y�M�*���F���ktv�a�~�h�}y�_!���'X��C�u�@?��/�7vP:��Q�J.c($���"%!��&��(9�yj/a��%�gt���4P�Λ/�,��1��q����G�wC��l���{H�p��!A��n�8��О��At��)�A�E�x���.V9�[Ⱦ�Xzۦ�t`C;BAOa>=�R?�{i�N}X�m=i3��8�j��(c��<wk{�kX�yjɫ�!"@x�S(�I�i��C��\�^0���k�a�b͏|��C���RZC�MnF	.�M�s�E��w��^��'cm�زQ54x%�4�x� }�	RBa��栨���_�EX)5���)�J���8��4*���M=��P}��׌,��mĭ�!%�q��"r$�o��?��z�O��sn���D�vԟ�6"��]��;��)"6�`;:Fg9 N�&n�Ҡb�bѠV�+���^{�f�9���wN�d�����M��n1%�j��G�����o��z��;�!��:ɘ��5�q�k��*�rŮh��8�b�FҊ�[#e�mn����9R��p[0Hqn��$L�nl�RP��V���)W�	˥EL1M��d���{Y�,Z#�rx܇�{�.���0^���`κʜ_W�]�닫�6O��~��Y E3��GU�1F�[gp*�c�r�,�0$|@L	�𔙁| a(q[|is;ZT�͗J�"�ġw�a�ӎ�,��@�R��P�4i�<��_U{U����N����hg& L8�k^6X�^��ǸT��.��PT\E�����b��E��M�:���=��nVi�����)v�V�֨�Syqcm��C��̍��0kIE8�p�EК/
@�۞�TE�t"����N�,�&	��������'-��K����
e���g�7�m�'��U�{�C�a3g�jTon~��<�ۮ�N�
����?& ���N�� B�m��Zݛ2uͱ��l�?��m��=���ZE�����&�s�݉���)����y���?��m=�4r]@��.� �`%�aY��3O"�|�G"�%�V�pI��;[D`m��|��ōf
��:.�K��W�Qm�i��f�����'1��W�`����u�
S�{}+�Q�־�,=�"���k��	 ��b/���Tm�P�]5�չ�<߱�u�$k�۷h)��fPI�Ie�M@��RZD=�o��<{ۦ���psD؃&�d>�ݠ!���UH=O��Qvj�b��m�5��7Ҵ����Oi~H��k��wp�V#�,�5�g���<��U6K�9]��;{i6�� *����Ă���tAM�o�s��~�Ԛ�0�D����GC�JF��ԅ�1��J��,��#�V�5�'OU�q�2�2��!kC̾O�[A7�"��x"�5��w�k|��J��X���М���̹���� �]�+���[>L�%���4�me��a:1����(	��A���h_s4�k��Aw�Z(��LT$��9 ��Tw�+�xgͦ1�2[x��T��1�b�hl��h�0��<�퀑�Mv��e�zmH=�D�M.��q�d���L.�Mw���7 �L�V6z�&8�&�
�
�a~!q�~����b4Y0�U&rY�'��A�/�9#����up�]�vk�����Z�y�ׅ���8� �30r�D��B�v8�Bl��{?�.`hl��P_,��}�=��OD�\�-n;�a��`g���sS]�~����5yX~?�w�P����GfP"�dA�Ұ��N���l���_�d�$2pp�®-(����H��;�����̈������VN=�=qɒ&�}�@F�?jz_�߲jO���xS��Ë �M��]���m���ҙv�_�_��pH���.뇶�І��-��)�B�-���<>$\b#N�;)Jyg�ގBNP$P�{�z6�D��
s-5��G�mˆG���b6|��X%<��7�|)皑5�Q\���O��%l61bTJ���D���&4ݸ���#�&����]�6��ֈ{�OIl�<J]X��6��ĵ��bх�<�s&W����^�� �T:�C��6.��p_�䣚���z�kb���a�W��
=�~�~�f�p��t]�T��?9%5��W�����8���TP>�L��wXՓw�_?���s-��zǹ����;U	U�<�XH��(�3���a��x��Â��`#������u/�Iv�r
�H�]�ǁ+�|��P��I��$�#�սsc��T�YmDo�����,�[4�j9,'��-�٪��vG�)��^����;+�{��%��<[ �������Mfr/��
bݧj	X��[���A��W��Z��{>!1�!�"'{Nk?>����W�+B,�U�ae��)�РU2���^N��.��PȄ�-j	�05ܛ2��b���i �?���5vHe�L�g����(t߄�rZ�iV�J�Ŧ*�g���\#�� @Bd��k��r�ן��k�_ӖS-��4��1Jy'\6��f��X��y�������ƀ�0A�,������Ӯl
�t���Xa��}=���8�)�DB�,��ŭ�ML?�9�![?��iu�"h�M9 ڕ�Rګ�1U���ol���f�qq�}��٥��-�E̍������s�"����6��~�i�m��|/��wG�sZvJ����������!~���X&'z��	`GQ���\]ա��ƈۚ�Z�t�C�M��LȀ�R.LI���x@eҧ؇fH[���(�4�D��gЄgv!IU|ХT��-։w
M�ƾ���Q0��]8 ���QE�t�^�Ɍ�X�و��$,���R�C��y�`���$N	/�MJ����<�N�в,ouQ ���Nv�� �C)���>IMD�ʹ�`��z��� ���BF�Y�ٌ�zV�R�U�WB���ȃ�d��_�	Y�'���ap�NW���aQ�����!�h�\Z_��I�>Ji)���朎R$������Z���,���vu	Ф2R�|*�zE	D+%��vvCJ&��	��r>3���}� �K�he��X��z9_d�HNZ���"ai��xoPF�n�-j���Q�T�n��E����IwS���7`��ż� j�0�0�/����l�������Ѱ���ѹ�F�A;ד��2�8X�Ǘ54b���a�D�*��` ��0Q���|�[wan��C����΋W'7�8�-���7K�J�k'�G���Y�����h��{u�niI+[Q-��3�9�0H5	7g��F�I��Gʁl�����un���(->!���5���&w:�}.9�]��DA:�@)�EF{�rݞЁ�;T��W�}4��n�}�ڃK�Y�`�t;E�
�~�����]OcJ+c��=.K^#M��&������S�����>�4yVHǷ/y���yl��ڲ�O�Xyf@��Zf��e-�ۏS�;p�ӿ5u��I�);~G����Ҫ�Y�~�IssUi�@SV��d^��bH9��ˆ��t�(1� 7���5xfg4{9������J��������s�Hej�z�����F�2�&��{�K����
*���5���~w���ʐj�f���"�Q���z��)�Z8@�A�X�J�ρK��~čc��5Db��,�������d�z�����C�8�ˤ{�;_�8i��rPj�A-��!}�!f����Fn�#
��f��'2�A�J�����:1�<�
�o8�1���}�\[�K p��%g6P���17Q'�}z�t�n1y{�ڏ9�ݹ��F_��h;��g�D�L�b�A�{+ָ�a(���q�i�!ܠ��Խz��j��s��q��H�\�%C�m�D��pa��3��d�M�S+w�mw� Qn�Fmq�ۦg�K(et<7J2��+�n�Fq'���v
��G4t�E��!T���Dv�2�����'[섀^t�}�nM��1k-�3ݨ�߬l��i�D��q֕��j������R����]��da'���(�7UYt1%!)��y�joM���M	�AF�-^�Tv��e��?�a�@]f�N�Q��O���RT�Qh#�ã����� �aL;��m��� `m^I=����p�?&�Ԝd�$�.�b���=1j�Z�]�h�&~��~cQ�q��3��y �! k�۠
�\=�/9���p�5ۧod�*$0���|�UHW\���p��Y�)}1١T2�F����
w}5Q��>z �,��*��ocP��1JL�S&�p>#n����L�J3��0�ۺ��za�����ɾ�ө��4�V_�i�oP�����m��S��C�k��\MEAҶ�ba�0�&�Zur���߭<㉲ ��y���ˑ#�z�Һ��@��d1�B;*�
�vt�JX+&�-]f�kӱ9��v6a<�XY��5�wW��X��`5���y�p�?�9����� n�����T~��1F��{+ �ǻ��L]��a��%��n����i��LfEgyt*��z��[
���&y�r���"�(��v�����u�#{�bk�_-�V�\IA<
�� k ��`1$���_0	S�_���sPZ�f�C�~��3(��Q���M<b��&[�M9�qԠ��9�_9�4�׀I6�ѶW"��3Qޗ���dΔvM�K�R�$z��	��RÑJ,�@��ƿ�C�K~"1� ��p������>n��0���L!�_'%����IX�i�ƥm��}׫��U�4���X �>T�g�}�y5��ʜ~����H��-i�M�(�,�&})b�	;��!��.�N����!Bm4K`�N\��zq�Jc�h=���Y�"��pIN>��e�H���(1��R��6~��v�iV8Ds�ި"��'֑�e��a�h��[���.��W�B�v)U��0�X�Pt���!I:�x�^�]��BC���eV��B9�T�t�j]L��u����K�݃��������y�3O	A���Qɘ����y�V�N+^:�?���eN�>���`Z#}Ik��ߣL䭍,��p%��Mب�a�]>W�y��@ǬF�E<��ݽc���	�ϒ^���l;(t�ű��f��	AaLSx�F=�Y�k�\��D���Z-�Ml��L2&s����1��2�ϟ�ve. %J\���Y6��M�	��!�vI0P�5&[�D�6�;f|��5'�@��+��	�Z|�g�Bn�S&�k�)�tZiƇx���u�'� ���WZ"t(�E|��m{�Vo棊�T�������nb-/��4v�r�_��#���߅X}�)�lsp-�w�/z�L�P��
��Gz���b� <h������D��U�/l�J`�#>�����j?�k�u���-�)c�`�����7��w�|�[m#��3f� 	���&���"H�K��0a�rH�7�`�C�_�mC���*ȊL��J���s�nf���KfQZ[:�<�<"�mR�7K*�ᐢ�g�׋�Y�&&���2d&��`�x0f�C;�*5��T)�8�����(/pl�0�?���_d\J���9Q��Ƃ�	�Q���)��(��q��#��[�@>�q�s��q�F�{���eŰ�����F�Қ��P89l���u��)���R�P:{0Y�j�/�O7�˳���T۬N�//X>���cE߉���D��7�IX��� �l̔<�T7��º�,�����62"�1�0{��q���2)/���g�]
p�9
��X�c.���8L�nO��B�E�|1���ā�X�����uM��Ǖ?K��p>�ci�`$�P���KN�����H�à���1���
h� ���ɩ�d�ў����r{0�b@�)�%2�.8���w�0O^i�Z�d+�ش{ge|vK��I��- ��а�O�/ժA�h����c#�D����{�}=���f/+{�U֥E�KR���U/ Bz��l�4%:�3���Q�_�I�9�DZod�Pkץ�c����iEB����"a��Ͻ�0	'����u�l��Uw�[�x��D�O@&|G�C�(�ofB<����}zSf�C��f�K�BD��w���V�ˊ�BhW�?�KjѦ'�	��_�6^�η�LSD��^h	s\���˦R���|�� �es"#�3�&@�ӿl����O����x�E-�O�ta)��M���5�A7N�:��Wyj������@��UR��(5��G���J��Nb@c0<Ĵ���s�>h�"ŉ:)@�q�C�\�?ˢ��R����K��^�8�a:�",Egy"�S�5�\>r�e�|Ÿ�rV�y�F�oUP:<��U3��� ����W�G�pt9����r쒘0@� �%|�ѣ^�������l锗��P�2��|�P�s{)=�5f�-Lŵ�fX�k�2H��`JG�P�{I�{n���*��%� ���p`#D��AM	^�����ռsX�A�.ڳt��x��eN����ln8���z1x�gh�݌�_Y���!�8�k7Jʘ�z������ ��e �8Ӹc����|���}G;��@zn�v~���N0L�,kԭ,'��D�b�mp�rD�c��dLwN�WwJ����>��}���`7TzԾ�H-ρ��A�9-�3���=��0������>��W��C��;�H��1�X<=��x	�,�,ƞ��|�$�H��c������!���OK�lYF-���%�T*@>���|��j��,w�� �V���%�|z�کe~cHW`����pq�Ա���)�>j�!�]C���5#�2:����fw~WC�z�!-z��&�HPU�O�u��I���ȗJ�3��^@�ږ#��YF6|���.����d�����|��z�4	�MT��[;]u7��P�q��jf�����M7����^�U�F^�0��h��`��8��5�\�����b�_����(�Z����$;V�J���b�ڕ�r�n�-��^�f�_��.M�l��F�Q�C����﷔��z�i�h2%�_���R����4�:�M�i�|_��^�LCa'�4j�hS��|�w���i��L-�k�D�%�l��Pۤ &�����
�:]��+��a�`Ɨ֖.��������6�T�[-gx��WT�~�l^����ã�XC��t�������rم:���������붬<��Z0�S��ਃe�HEC�e)j�Jb�>F�>D3/]>�R�����O8���44hk&�V�/!JQAIR�����7Φ7���k�r���іEG�ZB�Ze'Ԉ�����E"I�s��P���� ��݁�_&c᩸�A�2�˼p��M�t��ȃ� ����\�]�4�-�'Җޭ�@�����e<�0K���-Ȇ{f�.�H�y���ǥ�dH�)�;%F�{��#�����5Ix�gL�pr���[�9����`������$~�+.FӇ�!�_wޮ������]R�9�y��`���[� ��pD���}�`Q� �£b����EyuM��R@��pt�9%�g�|��	OZ��[��<��X��NC`�{�KiRw�b���WP/�S��_8�\����On�̓�4��� @�U�Q�d��$�T\�tW{�Z���j�Li�#ㄲw�RC2���9�~����îm���`�*�{�:И$}4�<����I�䩿�%ԍ�q,�ݮݾ���7�?e��ݹ�f	U�x�vCׇ~TN��NZ�W����%��/��^2������=�"����ү�4^��`�A1��4���7͌.�nv�t��Đ���w�G`����u��(�j8�O��=����Lu!Y����DR�x\4lM='|�-�̭��Ͱ�¡9h�'���6����I	�*��)�B����L�Sq���;�=wF.��bK؈"�:of�߈M�[������c=�x��M��)�BO������3�?�����Y�6:�t��\d�@nʶ��R�j�
�Lk�Pj4��N�]F��e���O�v��XG������}���F%�qa�F�˖ @� ��R5Xu�t
�7�=���OF7��SȽ�#�%#g��iw �.��n`Cv=ֽ�[:0�^a�ǈ�N�a|�"�eryp���������$��͊�tN��{�3�m��im1*�67NCG�~o�ϏgWڝ�K>3,�2W\�QF�qmy���t�rj�L��>,�y�U��p.S]-�2�_�_��:�����v�&��(	ӗ4�'������-} �����x�ȼd>$�UP���!�j�S��?��U�o�|���� r��C	#�̱������V=pڶr)%W��OO9��3��?ih�"Qn��v��=�%8��-hae��$X��$��6��=Ö~�,'�K����ܒ��C*���d#���|LN���hE�!��'n�Ak�T�?��'sJ��,��N��+C.�:t�� ��ܲ��=S��o,�R�ʖg���U�?h�R�ݣ�R�*�afX6�� lǜb�,�E�u�����-�t�qj㔘ԝC:"tTޖ����!���:q������7j�9LHS4���r�ԙ'���_'X �x��^�\��z"DA�W�v�eTnU�Ƈ���1��m�"Q�7ё�K���٘z52Nn���H"v{�żj�7i���טL�$O4����G\t}�H��N7�>eˡ�I�A
��䭣��BWq��K�1e`	Ev��M�<���E��$#�^V�A�XF�����H�F��j׸DEz8�*�����R�C�����_+]�KnɊ�!�2�WֻqY��q�P�o�u���k{�����],�������y.�D��]�#�v��Db�b�v��MI���5�)������2ʍ�|��tU��T,����*�YG��,�6P��Fse��X(6�u�����y�E���/�GeY����ť�w)�2��o~��Rj�.�{���L�[�w\�F{dkR�|z�P�<���)��G�ٺf���7�����w��LrlP��w�)9&�d*S�+-Xݪi�Ne�s��-�(\X�����3�t������?�����B{}��W�;"�+�Mqe��]Ut������r7��)�5=����?p��W�$K\�CaA��J�t��W��@�|��;�'���&�
(j�	ҵ#�r+<��ଢ���˶+�>�?Vck"��w�ۨ6-(�Y�x6�EuAP�R4<�$v�f(��ڵ&�sH{C�=�pߟ���H/��RSS��t�QDEE��J��~Π��^
���8����� ]��
�@��I��00%�l�I�Gi90�w�opF�G��A4�9�jE�o�A�̧�s��`�r��%�8�S6�Ly:��y���}|c�+�r}-����\���.:���D��~ i�,��aI"�Zz��x�Q��N>d��x�GO�ِ�%y��K�sH���P#6,8�(���_F�S.�=�[�G��?��h�a�{��&�^`?k�a	>U��.{<!���_E�@��±Y�A���e�*��������%�1�,Y�>�[ՕGʱ(s_�hc��,�PǛ��x�I���x05?1���LS��.x�X��x��m�R9���Vxÿ�.��f�BC���$`,Ss0���2C����y`�{c�:�BJ1�����m.�[��+����t���ϖ��xDBt���v���+T���
.+��#�\4��g�g�y�oz���1�~6+x
_i�����i�K����t�p�:2`«�F_>Lb��m �Z�/��N��i��:�t�,XQ6����f�w�î
Ξ
�C��&��_k/�"��#!�ݺg���Na��IcVZ���?I���m��,������0�T $gñ�����u7�ڂ��8�|�gь���%�H�71�"�%�#�m6�At����������оf7��u0��z0�	��%GĿ���jݯs��=.N+��$j$N��u�K�J=�)k� |��$�8�n�8�D���b�0=0)l�c��-�����b~�,墲��:�&�Qpư7Tf�g�P�1�ZN��r�A%e�����S "�֑Y�t�� !bmF�˥!ܷ�5x)j��f䯂JSH2�ȯYV�eMDp��j�p��d��!�ӥ��س%�����iNj4E
�X�����e����2l)�_��{��������Y9sq��}���)^�)�LJO0��.R^�����}���7_~<��'fɸ�����G|�.�W�p����,RNZJ�p9��4W��o�-38ɩ��1:���wߜ M*��Zjҟ�)�!�	M���ڕJ��ư	"�j)ӈ��\��1tt�h���STg��.l�S�vA�rE�_m�{�#mv}�:��E\�7�X9�$���nO�H�@���C�.�+���7�oi2�DZNߝ�7��� ���a�Wl��M�$����_'
'H��]�H@��	Te�s����x?��S��%��ņ�Z�&�E�Q�͐!6����|yH��y��K��=/��%0�:��vK���ئ	S���HCT�־�W��e��k; �m���JUu�>���p�ʛr�����Ws��RQ���>����\t�x��؆>2�Cc���Fv때2ɩm���y�C�#��]����x82�(���E�=���J�P���T�_^3�L�r������!�ƟG��L?��y�L�m�Z�pb�;�	�����n�p;a����K=	Ng��y>�aF�Y w��"n�-l��	5��q���^���c���b��.�X�B���d�� �3��L��cɫ]^�����������agM�i�Tf7Z���\����[ó�Is������3�(f&MM�5f� ���`]#���_S/��#>s��GǐҨ� z���W�;/+A���w��n�����9��ތ2n�3�37c)~�!�3v9˶##��>T p�4��Ty�C�|�^�s�`��r*��w{8�� �Ƣz)��G�
��@��U��G���Q�R���c��C2�2r�9��I\���=�Ѷ�+T�쳈��a<��)�GU���� ����.ͺY`9������c��d�S�t�f��1��A9`Xe;CC�1��.�9J�p~��dqy�żFlBu�i��VKÇ����ў|� ��%��k���rԬNʙ8�l��Q���͉��ʶ�Vd��k����¾��g�6n��ZW�v^��P�� i�|�ssԐ��vC_�ӯ5s?�tè��VE\D\.��!nhh\���f	���	�!��o�(E9��B�����J��Љ�th`�h���.T��s�A�`q^����?�� ���o�Ӽ7�P��E�P��pbL�v:�� �-.���9ˏ�t�=��|?x������vDl�u7�;!S/d���F�rf҄!�B��d�'yv�(ې�����5A�rhN�×2w�s�\V=^&�嚠F1�i�D3�Q�A55ǛCʨ�E,aSQB���k�8by��&�P�cX�R�<�&���Ȯ�n.�Y���%���2�D��)
�V�(���k#u��W{�#G�c�>v(G`c�0R��:iz\s�2����,��J&3������C`yq�g�11[t��Zr���{չ�Q��6�WH�K9�����m�Ό��� q"8�6o�I�y~ޫd�����DͲd��dS��WOX��l�9M����	k=,J6�uWfU���S�N~�-�ФxQ3�=y�J\u���7;}$���7�f'�Ѿ�J��I���cfs�����T�S��T(��⿽�Nk>�BquI�G"�]�U��^��3�H�����h-1����O]~p�S�2���
���6�=��"�]�O�;#я���� SǏ�m���=�vKs�k3��nm4����+N�J��}zO�!A�����n�o�8b;7t�)H��cr5�\�����0�m�^d�e%����@ʌ���	�&2��tm��W1H�u�@��z����t���E������{�Yᘃ�;r�7�ޭ�r�Ld�,��w��j2���Qy�V9CP�y
�Vj~�`A���t��܄�g)}	��D�+����P�\'Ф�{.@��x����q�m�`�%�]kG��OЏ<���9�~�k���i!��]#NA`Gd�P��f������4�q�Y?Q�	���i�����b����
�;�]�g��.��2�爒f��G"��KPlF�)1�{�{Ŷ��+��&3��sn���O"�:��L`�u�~����c,'�G-[UǄJ�?/Q^����`�SZ��i�n���&�Q�i4�gLo6^P��&��x�J�����3�"䮇�zpҟ�H�f�������]F�wX��#H� �k��g&=F��7�����ťj�/mBob`R��-���;��4�+��������o��` %h��=�~.������h�|Ɍ�흴0��'��1��,��5M�j1>)������+�U�/]��c���Y�Y`����qDD/�a�K�K�@�}���H�{1���0v�L�(��쐼�N�aTyGzرH`���8�8}*ۗ����0�VbR���:�h<sq�@��Fރ W�Ev�ށ��|���
~�h]�����Gq�]W�Y�CZ٭�~��#�dJSݦ#�o��!��|p���F@�)E���/I�.�;���%S���QĔ�Oe�Nޘ4�֒B�1�R�IQ�J�kN:�ҔU�,�ʨ����ٚ�e���w��K�҆�i�P�P#GH$���@K��نk��}n���6��1���0uU�x�H�cUG���W��F��ݻ~/�g�LvUv���޵���Z�=����O!B�)g��^{�(O'&����h~l��g!ZfDߍ�Ѩ��B*y���I���Vq��Ԓ�����FW�J��k��I�����T�5~}��~S:܅�%�+u��# FS
xsWRDY�47�˻H���eƵ�!���{� $& ����1��}����m��;�� ��T	D����̂a�WK8����k\p/ ������e���K	%���Q�-&�L�S��@�C�Z��w��;A2����c��Oq% ���)��W����7��)��Ӑ��
�)�Ȼo�_�ϯK'�	m&��d-�\�8?�'�?NNs�b}�K��q�j�J��UWH���xXه:���
Ī�FӃ5����H�K?C���/��G���޿Km˯���8����>�HT.�P�9,4@�hM�ٲW�A�D�����g9�x�0c���	Gg{Kæ�eCh�k(u�3�A�po d�Btt���V�?�#�,&x��P���C������f��K,۩�sXs̡���̂טӽ������.Xiql0^�a>/�(F[�#Z�l\\���r9�$VC�eAy�2m�y��O7�����r���y-�Pj�RǱ�&N_��(��"Q~ �]�Ǹw���R*�H�b@��a%�'^���ֻ=g�ȳ��fB)x�m�M� ��|=�cء)<�8�|�*���5�c����������)�6F�b���Wo��wFd���u���O����$u%�c�E��&#��l�\���,���Ƒ���}{Ïq؆Z��Ѳ�K"o�:�l��^��!����LT>}�F�(ԉ�|��I���#HW�H�75�j��v���"CY�a�8����њ&c'�+q��z��̌�$��k��:*W9"�;pM���;�cU=rb1m��BD];�a�!��v�9l26�wG55�3���dr1)�Ҏ��܎a�S�
H�щ�����-U_�=&�n�#�{9�����dw�?a��!5%�\/(�g���4�ƕD�f�vsB�Y�:_q��^n�9����4�vw渶{�s�&8�AX8y0{�Ō��Sp�5,�΍oГ:�l	O����������ޗ���u|Gx¢"���`�k���=�ɝ�`�9�#̪Y^�k�z96r5��9B*����{b��H���tho��K>h�ֱ*I3PM���n��*�P�6�{�!ͪ��J��>����%��X6�#��a�+^4U� ( ��|hE	*������|=[��'g������\����؁�p��(���M�̅�r�~��l�S����NRG���L�Ѩ�<���l�?)4l�$�F�HH�76%�'Tiϝ�"��+��ڱڥ��,b��4N?�/���a"��z=h~�PM�,�N3�1=ȮA��uyuL(8�J!:�3C0�aξ+q4�Q�8$��0�L�aE�}�{���0q���^oQ�=vG:�ȓ�����TU�fb���邱J����_���'�kK!��z�{�6/%� �+������`D>���]��M3�,{�0%����>j��!��"����a	*�}��t����bl'�A�l�?�b�T&`b+ՋV�"Yn�o����b\r%�D#�]�ܐ�ג�4��.*:�؉m�����*� 4h�1?'C���Ʌ6�`M��d0a:Т)C�g��F����.r�@%3l�������,x�\�EW-C������o��8j��K�Ȼ�c���Q��ߞglU�I[su�J/"�Ey�0�<��l	Mt&8��/��
�����ܠ�=f����ޯX�k;K��F�_I1Hxk��е��#e�1�,�{�W��~	y��F�/��l0��q�7�Q\��W�������|Q<p(��"	z�w�ʵ�����'7"�t�%�	=�1�������A*���fJSzoUAT�v�@�ƣ����Y�K$Mh����f�A�V����� w�h�?��Ø'�Ǵ����6�v��m�qju	�����a�G���)��vz���i,�}�����;�8�a���5�5���O�%.`������!��>(�P��&~��T9a� ��歒�խԯ��xOzZ��4ۨCTz���	x�HX�[z!�J������Ҹ��Js����3j�����EV�~��d��V[Y�zc�^�Ϝ2�굌!Wv�n�D�F�#�[��J0�|��.��_f=��rj��G<��x��8�G�"�b��ո������L��S񦺲��=3�-���}z�����X��1�]������@C�ym��$�~�stw�LT*:ޑ�� ���W���*nԖ~FuCe)L3�q�I$*2����M��N���Q4;�pY~�Ƶ���c���=��y���rn�)��Z3�f�)2�]�=�^�Yk��n�ƂܒS�	Á:O���Afcd�гZ��)F�Ğ�3=�-8@F����f���1.d�W��<�`c��kmC��}�Nm�Cz�jD�e�RZΚ�ј��?7�����<�m�dU]λb�����)��v�b�bLT��bm���v�	!<x�p=��,FV�e�L��,�-��46���{x^~�(��b�wJ�����j�V3T@<xt��:����4�xf�S�sKڼR���7v�uC�LiM�mFE�Tk��aҦ	���pUí��Y���W��㧿��Z��#X��a_�-8��{�M���� �3�"ՠ^��0����]�?x�>����/�����`�C�r�D�sげN�4D�R���@a�\�J}G�y�p�{#���g/a���O�����N)
���y��=�f�܌��/������}��b�F
�:����Y�l�
&�9��N0���)�)`*�����Tׄ��qK���ռ�7�����bi�W)�;�eq�]�ۈ`��uAΞ^[.?��OK�Zs�톇�������H�Y�\�����h����9/Q����8�l٣�Ԇ Cvl����K���,C�5.5�-�h��ks��G��=s�g�	��x'��~�b��~�@�d?!�S��w��4t����ԃc �W�c����g~�"[!���� a�(���_Ҏ�,�h����=3����%D��u� T4��"�2�.�D���}Z<�!�K
m�8Ā�,�̖Z���c0i��Ny�nDf����v�xt�KE�
�z�[WB#��]b�_D{c�hSx��-��/T��-R[���
ʂ�^��Og��F34�����ؼ��x�X��K6)�5kt������3o9��G�`�n�IO�(y�R�h� 6�L,Gu�S�7�@D/�0Iý�eY>9����y��뿭u%��ח�ݾ�^���7	B����2�ѝ��s�$���[}��΅��
`�MƊ��7�����q��K��7�I	t�g��{���q��U�:_��\	����,��E'{�[�G$�k�#g��WJ�vo��1�;�� ��M�6Z�b��_2Q'��x�%9��ܻ$6r���)m;�a�����izBX��N���%�~Q��ʻ���k�J������F�}���w�/�ְ=<͆Xy�!0���t�Vպ]Ԣ�EDQ�S�>�������ɸE\\S�z���_+�u��y�8���=�O���>3^�oY�6�L�|}"�l�6*�����A4"U�.Y`�e�>5�;�u�xaOT����7)t�K�ʬ�Z�n���@~t"%l��#�nT�-�<�IEW3��m*���4��/ 9S"�R��:
��6uIe���k�.�}����j+KN�"y�S&��No\1P��:��yόF��l�p��J��ޅi!��qzB�*�W�{���&��֌�ܲt���,���C[���Z_<$����~� oi	P?K���k��l�k��\O����5�D� ��,}�;L0����E�.�
vjw����:-mKs����c-���Ά�%T-{|��@�/��?�q��U,��;ܘV�h��0W�������М��@tu4.�VE�_�Y�����ܳ�7 ����N��4���>A�T�s��b�؎�9�kM4K�5���O:���p,����ؼ�9��!1Ƞd�*5EL��{@9�J�8�wz|�HUA0��8���>�7(&n`���`���~�B[9oE���m�ҒGbU%�A"��H׷��Q�BsG/�[�剭҅T�i ����l�H+M���s��j�z{����3�v�	=v��z̘��U�Z��1�#��^��3,=��=�	�E3�ztH�%w�]4�vޅ�%#r9wX�����]���[` �LБ�E�����:w���]�Q0���FF{\[7Ѻ�s+��x�#��OT}��;���|s�@y0��ǥi�O�4��n��VJ���y�!;T�L0.��*q-��y�|,hXå_;̛��N���̠y&(�3z_�R�4���6�4��M؂Lm�)9�A%�%���e��.mk$<sZ�$�"߇cm���|�_2\N�0��Ȋ:�V��֕�RE���1�N(�c�&�<��{�f�([b�C�&�@��xY�q��2O:e�ph�`$�Q�[�����~t�[���j~������w�r��G�x2NS,,_Q�']t�iD�� � �i��ɸz��f唬Ԗ�қn-�Sg�{����y�S�ns�qPܳ��>J�-���E�V6���݁��p�❽������H��_���i��'��x$�I��$6�@6���y'ͽO�8vn�����~7H�X%0gN4����C��^v�-��¤ ��4ZJ6H���%��՛���kw[9�\9�0�.z��P���d�c�MO�r��MeM�?4��=m�.��BZF�{[�͍=�S�v��z-����~��)���ٗ8�Mg�/�7_�u��P��`}�n�:(9���X#ʤ���a�u=��W�4���N����@�A�Zkؚ���dA��'��ݣa���@��p��xH,+LF�^���O�A�x'�"�#��\=�Z�r�^�������ʺ6�<O|���Xa��U��F�(}��c�8��=n�3��<'�^-)@ߋ�:�u�Kw�:�28	�V�$HG��d^��J��Z���el<Vi8����#����72�e0�4�qe���.�b4��T*���sP�"0�EŃ����~T<��n��������&կ�4u��$��n"W��v����O{�2L|��ktܳ�y:*y@�q������*l��a�<3!�y�aY��:)�����;�ԧ��	���T���XvL7QP�C�,�ƌt�_$S2�c,V���=+ݶo>����˺�S�z�U{���}3X.T}�p��|�0;���C}~S���;\f\����+�W�����RS�R,n��?��0 z"�U��'5[ww�����r�D�
���;�e��*-F��5�����^a�+�����Gԕ	����a��A{n�i��WL�Nz�����nj'>�� �nr�o�������$����sNYs\�A�(� \w��ՉU���W�UM��0���U:��mR�5���P �AyX�W�=玙0���&��s����h���i ��o�.5�����#E+�[�"
���K��0v{H�E������o����t���T�dq��]�:��-a��BʀͺF~Ƙ3�;�����Eܛ���|#xq��<]��B���Ԋ�@�)�������;�Wv���]���ҫe�qkWy-j��P}��y~�q:��V~�'E���G��=���MI�4�Q��V�I���Tc]�}aG�R֑<��������aƙ�:6Y��	�ۄnq|��1�SZN��/��aƖ�3�a�F�pk��Z3-�Y��)w���+}���SO�+!U!��mý���V�]��	���tb8Q3�	�� %���Asa��c5˘�e&}Cm�)��0y���b	j�7�dT2���'joסQ�?NޡDܴ��PG-� �L�Ί��gBC�!-K%��l|�m���%�[��)iɓ����dB�������E�"���B^�'h"�}�C�-|�/z�P�J�7C]%�0��?��<lO)�/``�i����<��;WB����\'�x`��ሰF�����Н+þ����?��)*�9%P�Xx۝�l���b� BZ>�>S��&p��M�=TN�qb)ר7�l�I����ׄ-p�s�4���^{�#j^��Zc	���MT�.~��O�)?Ԗ�)�v7��C!]s������9H�sf-��,���ޙ.�7����٢��"u8���C�]���������b����~.F���h49��eb^�gt[�3o��:�+ \��XKY�c���d����������Z8Hɱ�h$�� ����G�U⑙��,zv⪮����(��&G�[�)��gLz��f�b�����3y�w�\�j�O0H�X�٫��S�H�#��ɛ#�F��m4"�۝4�v�U��X�ѥ9�v S;@4�o������i��/���K��[�Ҏ&�QXe@�Э��^���r�-ŎZ�������΃f��;��U�E�Y�Tҝ��Y�ZBG�X�~�*�]1���X��F{u�y�/ͥ�,T���׎����Ҁ���d��5�JN�h�zm��P4<K�M�e�0G�6�*�`@�A�6��^��N	u!�٭�h��j'L��.|7ЏU��s:�^�C�2^׶sߧVTS���� �S�8	߭�ą�,D i\�7�2�MJ���gi,XU�cH�.ҵ�	)4S�=�]#����� P4<�*C]ҵ�4x_8ӭ�+Ife7�w�cG�gud˘0�z)A���'�y$�zD},9�� �*�XQVJ��vJ��HF�43'�0��a������F]����DQ,����}G&=
ﵤ��z��nG�� c�v��'�'�8���8g������؁g�w�\:Mi�^w ş���+xSa���C��]��r���C�}���?�E��՛Q7��45���k��V��T;(��G^������Ⱦ��9���L ��hk/Dkq��:%H�@�-:��k.pe}�:Z � ���=��$�)�+�b��V��}U�V��qG�򬎽#��Ù*��}��Ƃ��v�lL�8�愙�yխ��l Ā�c�o����� _N:$�C�{�<N��o�|>|)�x)YM��=Pp���������-�Fc���!I��r�:�u0trܯOHZ����o..�z��#�0\��x�\�S���N!}yV���������9�ƅ�|%I!��]�B̓L�p<7a��Ʃ��C?���<��5U@����e�5< D�>c}y�Zx�S��!�ԊDtb|����t@����Ǯhz�h�2��i�T�;w9�Cr�1)����]6������*�:���V��T�Z}��p�L�h�D���ASHRM�
��o6І�etӢ���OVO�Δ#��oF���9wخ�!�m����q���	�;4'�$��o�y�8W���ٹ�����Ux|����<4��mw��$��8�����X!P�t�������rq���䃲����vɌ1EY�����e�{_\)l�`��֣�S���.Kޮ�$Ȳ&�nP,�U0׎��������PG�c��B�����c}G?9��:�_���$y�34�b�9ˀ���OU�-�R50�Y���ꑔ;�BCnC����V O>W����W�&�����@o�;�a��+���$z/�G�Ws;����07[|�ϥ� �@ulJ�M$'u)h�W�#$W(\<��
y�l�ݹR;�"��5�����4Rx�~t���������6��S���b_��1��=}�����^2]-N���>���.�M�gFy!�}��N��hM��d~�A���4he�r�Z�(�uE��K��Hzܣ^l=ս�;�\>�@�p����)��h�L����UYVN��,E���m��Hl�p�'��5�C)jj��(m�am:n>�����ɡou��4�ꟸ?/�|]�֔C&|�6�V�-'�Տ���б�1o����z:mY20�0���(TACQ'c	����z'�יp�u}�.*��9�9��_`x�����-P�ZऌDr�N��t����"[='�塒�|ά�_�`��m&��!�1}������5�2�Y�j���7�����C��`+S��0��O��I��w��sO�4=��;�xm����"� n$c�d(P.h��F6��Q��a\]F'h2vK�w�+�lf�G�J�,_@R��K��< lj<��㉿�k%����=���m�2nT�*Y��Z|��f��)�mm�
դi^y^:謀Y؏O�|��gP,$�~�&�i�*s 6l�6�;�����r���Xܰ���e1i��i�2l[��$ǆ��:��ks��Ɏc�W�md�ops����_���P�^��W�B�>f�E�e?<�*�� �j�x/~�L�ɻtf��lu�r&��CCP�h
_��o+��'�2������x����x_%�R$��?H���R�*z���:mz�m��j����|�`�Q�6bo�q�	|F��8�@"�G�(̝�PE1�։���!g��l��W��U����o��>�7��.��}����:&�A�k�ŵ�e�D�vL���m�fS�W�rх�>�6g�*)��d��!��;�ˆ�VmX�;���ڕr���8;wy4�3�D|���X�Q����(��sai�s�˿��1���u��B<I )hUw�'��[y#}��ez���h���p�=��U��6�(罎ɇ[ S e1���,����)��7�j$O� #j�8i���%�d�����/�1�C� y�<�z�[[�['��]�������v��k�t���1+{����������60�g�*����}��*R�<�����EPNS�@��Z:�z��jE񞃜���t~�E��H�m5?V��$P3��T��k,��2o����ú�j��M3��>��N��ө�2H�s�L������]Qȣ/��!����*���Jy��'?~B2/A"C�Cg���p�dj����'dWb�����dp_�H_F��qH�5�/ec�p+�T��R~�/<��v7�T��'_�X�ҵ�p�+]�kD��W;m}Ciڑ��F��4�0�\9���#MK��c4���:Q�I��C�t(�c��|�[����-Hf��͗��� 4�*�̿1���i"��Ư�	��F�I�rH:iqv7�OƔ����Ս1݁otJ��e�.g��@/|um�<m�jŽ?�E�?̈!f
�$�����X_������U��l�ߞ��j�`�=��e���������q�by\""�����[s�}-�1��S����5�A�Ō�;��C�uW3�9����$�
�*M_��]�7�ʥ"�"� �Td:�GO�#�qF���9���C^0���o�Eq���h=��&d�ipɣ4mپ��ҹ�?ćהpU�(ۦ��ܦ�YL�x��Q�|��m�xq�o��Z|:��	;Ps$E*��'���j;�������X&�eq2J�[��/gQ�d'�W͜]N"Y��UYz�բ�� ����v�g��ǎ�ƞڳ���S�Ȯ��TmKu��_���g�}�?�V7d�ز��P=Ue	�E�"N���5��i�]S0�o(|W���tT�a���4O�U�iBx(��Q��F�0�жw����}�D�*��,��J���x4[�k�S��Ǧ_�t&��8�P��\���MW� +�!V�M1�-?�S�$ ͣeޙ���f.˰uaiZ�d	��E8�'�
���I5��(�ؐ���}�?�a������=%�&4��4Ө
��1�?���B�܀���;c��N���tx1&R�̒�5_,��)�Sy־/���(*3�ڶ����&e�c�>�j]��gA�`V�jzҜv*Iح��jK(R~g�������3�Z`%�7ke�uG�@�6z��p�M?��2����
e�~�O$S�觢;�>�\b�_WU�p�d����ߝVX�D�T�:��x�55 U�4�����(����ya���J�b6W�AR흰���ћ=��snD���n~0��"h�(M~"��4��N��*y��,+�?ɞ�ǋ>e�ģ �z��;z!��Ypg�|���	j��fN|%�B�	ӥ�Z"X�w��~9�uf6�0�N��5Z�� Aa�\�������$�ĢL��N�ݺٝ[�Co9��[�8Wh.�~�<�݉�ں:�"'Ov��},QD:��ƃ.��!�L�`*�x��.⇿�f=�m;S��VK���v�J��,��
a�e�m�q���Q�;��/���b��6>�m�`��`٢��G3��≸���[S�Ƙ��7Ŋ�(�������u��U]�Hӯ�x��k�،Qr#�}�>@�c�+�Mz�z�߈|�׮��ˁ��.�@��{a1�5�hL��7k�_�e�ֽֆ��ϯ94g��v�nR��ԡ��^�&cT�9ŉ��ms��C���<�8��?�1�r_�	�5�[x{.O����\f\U��	t�5w��I��~���j�#�����s��}�K���QEc@��T��]�݈5����jV�;b�Η.��-ݭ����FRG�J	x=:��������Nw1�U�l�����Y�<��	��8/]Z�-��Ҕ���0Z�ŀ�ꥉ�ְX�Dm7֯t����z�H�{naX3�u_l��%��g3H V<�W�#ȒWG��~��`lϡ�I���KV���g7��x�Ť�����pК��5�D�	�"[H�����NH ��J���{u��"��\���ǲA�y��9�s`t�B��@w�/p�}C$g/)�s����r(��qb5�|����� [�r!=�G{:��3�������7�fx�,ǸO���ǽ]G��_߈O��8�mJ�2�K��e�:���A1D�a�_?��x4���hߤa8��v}+S�Cyu�0.}:����xT~�4d\�!�6[V�ؕ��q�t��yc!�3����ܿ6|T�l.��Z�[��Ao�L 2��sX�(�r[Y�^9�L�Z��Kw<��q8?C.�m��s˲ı���\�V�0��[�%:]�?��됳�c��(o�;ʘ�����b�lb'�\M~ɭd�����R��8:��Dr+�QHT	I��z��Kb��#3w���<�?D���Ti�~�ᄞ�Z�ۮT=/���I]��o�!7h�p��v6�`A0Ҋ�8���� �g}��E�r���t6���#s�}]c�?Z�im�iÚ��?R���]{1'x*K}�ڭ�2h�<l�i��Hظ~��.���E��y��Υ�FC*h��%v�m��}��̘�	��۴%��Z�7���/��)���)�ķs< �Uh��.�G��Cv2���蝥n?�wfiM�)V=k�@ݧ/�N���ZG�<���Q�ǜ������7�ϻl{������[]���xaZ�6��/��_[�*V�� (��,[�ʀ!�KLf�r���ʡ�F�I(s[a\�6D�7�u�-����?Nvi���ĭ�k��7!QG����;D� ��J��lsLy�ȍWG���]=2Eb�(����
ؕ�Ñ���B�0��w���Us<�����.�9ڒ��a�3�E=p{�E�mk8!�]v�C�Qq��$��m����e[Д�:^��x���m;�6��{1ؽu���+Pu�fbr���}`׬�M� #b�e�0��2{,���BSBءԂ�kz���;�g�����5y�c3���<C��\�썒7ΨE@J.�u��>�aL�J��.�'p�)R�:jM�&�Y3�%��JS��ܧ�M����c@�,<�n
�)��Vg$J=*��c�W��Ș�J��wA�}��<%���5�6����	�܍_�;�	�?��/��nh[�h�\�+���J+l!�*�3����M��B�G`կ�>��ЍQ��.v�g��-[$�  ?Ō�ay���8cW�{A���j��B��pǜ v�`�E!A�����1��i���u�87F".{�u<�9�܇��c��-&J�x�R�N#O�f�����=v�Y�v]��gM��1������!_ء/�ɋ
�� ;�!d���s��N�Z֟�aW49�O|�j�ю7�z��<i�,<��7��]I[��D�s"�\<Z��t�>t�&#�I�EwSj{�2����m��	�Ai�(�3��u�`�C%��Ji�F���<��i�+7OH����a�푯��$�#G�Ϊ��kDwy�U�&�rv�`P�#ቨ-V��4fu�����M�{��Mo�V�u�2��>�^V�`�%�W�<juq�	�I�W%��̖oyhM�$�S���F�δ���,��ݵklX9�c[2��pT	X�J!�T߃�Ol�깵��Y[�W�u�"!�S���S8e*�s���+#)��٬7����L�)���2��΂)[j#����D7+���m8�����r�Ui(��۩�~G|�I!�Ǚ
:ܚ��fc�U�s�dT,��-������0�����S���J�k�o���u�"]Z�ʣi��[fgUUچ�%)������;`m�ѕ��\��f�|�Zy.'J��nNѢ��0A��%�){H�*�F����a=�ݔv*�cO�]wNI$V>��R��-�7e��Sk��?&�:��	�kج�
}�g6m���5���(ڔ�C�mr�3ޠ��OZ�4=_�)5$�#O7���/$Z���t茖��X��'��:�@�ʱ��(�:�#�?
�LU	��(��RZ�8�CAr���`�`%�Τ �/=��\�1t]�H���Ԝ�3��_�e]{��7	������K�rnJ�wbW��(8��uq�N�9��l?�`�Y�����E�tKp��{y�H�����6 ;�Ay��ڀ4��*���sYZ@6e'uP��z<�^����A8r0P�,��ŐM��>�G��p��p����oMO��;\���3X�.��=�@T/�Cm��kQ����F��� º���'Q��0��n�|�b��T�������w�W��W!��Eޱ�z��0W�d�V��ـ��ӄC&m�Gl�(�j��ϝK ��\V���-%5qJ&B02����z(i>,o���l ���O������ґ�_	��C� �8�S�^�q=	������t�SG�	����A�P�k�V�70 =�qks�AZ�,��9.�����H��k( ��|v02�)�^���;��o�k̇�:�I��b��ϓ��9�  ��w@F��rN�P-�l�`��8�j��}�G P��B���H:�{�G~7�y*�T��SLoC����I+H����zk����}�$8*t�S4؀�D��ފ�	���$t�`tÝ�!P��<�<OY���JP������Y��C��bЛR�Z+I�r�a�܁�� ;j/ ��3���"����6Z��(I��>'�I���2�g�3=_0�jP+j�~��%V[�w>'�\U ݫ�Ф�pQ����oͳhU�2��1��><i�B� P��]e	��>Z�*,��h��|Lu��l+g�7��s#k~f���2r-H�,�VB�h]K��#��m���ү�)	�6���\Ϧ��dt&w&��t�]��!�#�K�h��e+���N��=k�)'��ޣS�&�xb��A�L�w�))F�.���S1���lV�3w����nBXܤ~7�,H��(C�t7)?P��Ω�H����a�r��>	�˦�?��_S�[1��:Vi�&������\���[��n��te[;�\*�-�k.�}L�l��4f��6�T�
�!�W��ܚ_\!%�j����C!	�來"�e\���)+[O%b >�_p��K 0���7���,����� �)"}/_+�kU�U1��sw��
���R������u]���GX��g�Q�O�ָ�[��t{�&
e���Ԇ���E3pU[d�@��Z4�x��tN�.��u���_�F�&F5�Ӈ���`��e��Q��Xz�Y�����l?h��A������ׇk�
D�&\2_�U"!#[~�V
C1�l��Z�Gro�݅3�;V�.���}���3X��_8�t�g���}����V~� 
�w{8�Fn��%���q��*��z���~P��p��/�Iv��CuP���e<�����$�#_xJ}@���ti����>}t��pϘ�_��{��D琰4�$i3�Id~�a_g���L����:\��8�e�E/���9$�/���ī���u]�$���J &��t�ӆ.��vY�a��9Ds�$�ހP32G?9t�[+��,��%DÝ�S~�J��0~��)�"�<�S&��&�> ��	��@�Y8*4:�%o�0Y�9H�)9�ڽ����V7}�o�@�e��t3b؊���9³�����Q�͏��ĵx�h07��(�#0�r��௣|�t�������.�"`r�H�6h��	�at|>����5��b�(@P`ţ�t/"�S0c_��7~���E�t��@��%voG�ƒ��>��)�_�"����a�`-���qǮU�gN�'�=�kpk�!D%�k$��٭E>+y$��"�)U�
ݥ��)>��S�L���=�u�OJ�VX,��;{�^��h"��x�npLM2?�'��rO���`����c��yi)Jpד��U�[n�㿯�l�����F_6����Vžm4��ɜ���e��8� Pz��*��f?�k�~�I��N�@ ;)(p�r��Mͅ�l��v�VP(��	�@0w���@�,.͇T�ͳ�fj�fȴ�� ���J{:NK�M B-�y��4��W@9o��l����r}&����n���w�g-���pPM�~,?�;Њ�4��5�ʨ�|�J�ڦW�g�[^�F1D�&�5Ʈ�|�
�UԩH�4���l�6�51mĬ1����g<X*�(7E �
a��;|�/Ԉh+��ȅ�􍄨��t�?�/`�<�ɟ�-Tۮ�#@ʆ���WP���	[��'N�O!�Z��á�\�j����S��#$�E4���S1�t��'�Hb��K8���L�?W!K�*��P�8����0�$� ^�aџ��%��mL�o��իn^���'���tz�NP�1B�}ek��#���Y��7�~�u�pc����y2�KR( �oh
��_z�dN�R~�c?����]5[~|��;�91T�9��>j:Fa3���V��T?Ir�09�e�]���/lB"��{Q�W$�͠�HU�|�c'΢�bݨ;��Lkezn} ]oF�?`�.qΒ/�ff&[_`ے�-
�a����_���=,o����r�`K :XV�E�4G�@J����#����wŃ�>A3~?��-a�(�}����j:Ow>�`�c�:Δ��z9N�Лn}X�����frMwt�v�?kٮ7sx����,<m�]މ�$u��	G7`K��j_�	�-���e��hzk&~�"ɰ��C{2�(:'t����:�������U"��Y>D}R|լ�%hYB��##��=	IJ�h@�i��_��|�/�*���ލ�c8w� ���{3TRhk��w���f��ל���uQ`��sY���������H���/�sp�D��0sh�q��G2$>`V1�G���	̑G��pg���WV/�d��aFq�'���S~zRc#Y']�;W��k�ٞpf� r��~����	W��C�J��k�\M�� |~
���0���ݰ��_ʊ�����D���<_��h'�`�-������7����@�
�gGx7;�VH�(�9D�u�vg-�S�ѥ���8<�y��)bX�G��i����`_���8���������u9����Ww�q��ݰ/T���*��v�'V4!����h��*��P��-&|y}VcD�_�0,��{,\�9��4���@�L�8xVOx��Q MVQ ��x(��{���_M�D�5d�Hջ�vR�^.e~�[���Pq�7 ��de{_�OԄ���xU����ػ�I,�C�hBcI�.���XP�fs~��qNQ^�x�2S�J�#u��tu�_% 6R�{��&d�����vA���|QE�&�z����#�+c��+ng��(��Ĭ�(�V��T�,5:����sȵ±���e�;�������H<c)���iq�g��~���������OR�'m�u��D���$�����[Fox��#`�)�.ܕ^�Y��t��|��a�0Z��:l����y�V��\��u7�̶�=A�K�!��/�=�x��;H8f�Ѿ �a�܍�Z�(N\�}3?��G	�0U��[fuΣ�`|7
U�ͣ�b��$�<�E�t��}�5�K�I���W�x�=v�%H������i�+K;*�@)�na��V�t�挺��h�x��G����t�f���3�������%H�B����&�K�꣊����]6�����g��\EǞ#R�'�m�������S�#��ĳdf����q�Dw�E˳@j�?��0�|!y��L@��A��X
tn%#Ɵ��$�p1"1��q����w��m;ĊH?��.	�%Ҷ2B�qR4Z��Ch��IN�L�O��૶�z���7�Q��vBO��꾼�ʋ�B�pݎs^�4�S&A���]0%�c�1�6����?��f��V���<�qYy�����W
�0E�"�N�AFL�Dш�l�?�@�A[?/�`/r]��Xi�I�d�xtA곤�vf��n�� ��N��g��6SQ�I���/ �.�"F&'J��0AK~-��j���\x����P���F}�������_���0�D�}j�}J�;�o���BC��#d�-���Ϸ|6�8��~���y~(�b�S�Ee4��GLޡ�\��Jr���'ƞT�j�"��;kiF�y�pF���S�v,W��,?�����<�:`LJ���a]�4�mn�����~(b��6c-۔0�����ު�N�.�������?q�Go:H��v���a��ۛ�<C�ֱ�^7�� �Ϟk��7�c��B=����B�-�Ggϳ�e#�")b���d��]�<Q���
!�l�k���gB�N��V���/� ����-���2���kO�,�f����͂L���:/y�) 6W�����Y�t���T,D 8��o����+{ئ�e�����c�<]�K�s:���>���`?"W��?���c��]�+E{�44�д!���H�U]%�or�:h� ����{ȟ/+���7��;��!��qzk�8�z�}ﺎ������n��6Qo\��
xR���� �]����!CG�E��<��@7Ei��}.�,��y3����t����*��.u��E ����o$�=�8N�q��J(��w��at$�(��s��������dJ�xy�(�cn�"�q8Q���H`�6_�D��biD�����C�
�.�� �RD�Q,�|(bkB�(,JJ�����jsN��z���R��Fa�I�p\`�M9VC���y3���� @���\Y������|�9�6���`,�.b�Y��=�5FwV����`�I>�)����ޓ7�p������S�����w؋Wo?H\�.F�r�߲gM�m�uVl�᧻���P�	�0̰�D{�9,�6�|�rڬ�y#�v/+���F�	y>|*���"�u
G�dΣW���Y���D�׍ώtKB�I���I�!�O�뒭],�*�X�����V��?�o�9�\�*��C��t�҃t¸�ԡ��9���˨���b=�h0�}� �;�۴��y2u����k�z�cO&�ILaҰAS	�獣F1�?��R�h:[&>�
�ͦ�V�pe]�C$틽�P'�t�5p#�M��Y���gEӴ�N{Pc��/�̕�.�W�+�UY��l��l�$pg{x]��s:/�+�0���-��:~'Yp�t�5\!D�\v���lP���)�YQ�	��b�c=��"����+ZNK�=<�J�hl�h��Ũ�#Y� 
��w�Ǧ;���޴`¿�g1�<~���?s�̈́�ytbU�qh��<�6oa����L�e�_ˏV\���oXu�l�a�U;EZ�`���}���e
��E�5�7;��\��$]0�y�@:�\~��j'�v0���Jł�2?��,�$����(ܑ�J�c�����OAD�$�+{ڷe�^P >���F��;����^@�3X��P��e��Θ��}3SȬ��e �:�ĵ��w����	�����w�@zns�^�X���Z,N��HG�Ap�CI�//n�DԎ��Embͽ;��ΧQ��ͱ�ݫ��°�����r����gWX�oJZ�N��i1�6��t�V#d�O#���.�f�2���A�=���^LƳ���C���*&�[f��y<c䯳�C�C �k��i��94�1��^G"���f-��` ����Ea���wa>9�O��*)D�4�%L�³�@�H�����D��-r�z���z}�H�k��m���E��:����pL�\.�����窧-�W-�E���mb��}A)����� �a>����&��y�v��|���!��M<4G����Oŗ9�M�֣gK�(ˎѺ]���F#XP}\�;���wy��rN��_)�����M�O�-�v�U��(�K�`z~�P#䒨��dH�{+DZҮn��>��د��D�0�UfGrZa|��|��pƲ���)�眍PgDQ  �2$r,V~'�Кn�d��U�z�!sv�|���Q��3R,�@��y�R>�������k醺i�s��0�*�n ���X.���WQ�n��5vu����KZͮ*(�c��Q���
5�R��C&�,�t��F}X��)`�q������`6��O2MG���7�`B��S�I�{w�s�߮?w6Y����<����ڰF#���x��`�2�DC���j�'�V��>�]X��Ń�T��%�FL:�@zk1>C]�8�#�^#���a���O����S�v.����czX���"c��:�q�yC������
/�.��Z���8ƚUua,u���%�nÐ��n+�<��]DZp���(���i��DJ��5}aS�<�2�k�e���،�(��[Kj� g�j�Lr��KL��w2^�y���k��F�R���R?*�W����ր��XS��%"}w�7K܌'f}j1f�������a��W�b0�OC��7r~Q���J�Jah�f���������e��"k:��1wwZ��j�]#�{&ir�\��T����H�ug��=SN�w�o� ��0�w��W{����q�EA"ȧ����l� ��D]QŦ{ZA�<�Mc�!4��j�����SR���n7��
�*��Vg4ac<C�g&Px��*�W�u��%���\�;��t0�*��2�EhDux�{��rWH�����|�96S$����O�a~ŎHn	GM�i�`Z��v*)����!F�A��nt
'6�y*l�{`��5��$����b�g��(/4�v��S���p�	 �
Vg @Ya*Ұ��)�|?���rޛ������s�I'�b���zt ��S:���f!p��~�f60�=�J`jo# �~���������7��8	�Oϡ�m�]wQ�[Ow҅>nѴ���4��;/�Q*��R�-p�v�$�4�R��Ћ1��e�C#��<������fI�#�Y2B=L�lb	5"}k��+�*�ݍ��b��H��9���ϯt�Gz�y#'�#��1g��JNI����%��4��N���ߝ.�d��E�H�&n�}��/��,��*^��G������)���3�J�2),�f~UE�bKz�>�1�}���_��Jsj=���T=��H5S��ׂU]��4m�L��� !)h޻�w����&^�N�R�M�lK����T��(�?��`�v�������vŌ�%� |>˃�8�}#��f
��
�"U�?� ������M�p�r���y���Ei����� ��p�Ɔ�Z�2&�#0�P�J~�{4���b�kGP�ޥj0��@
��Q�8#�*�H%��d�A˖ܻ��ũ�hr�n�#���1I����$�+\M�N{��2n�=N��P�Wb�+3�i(�=f������0��#xZ����`��d��G��Tƅ�k~t�����U}���k��+���R��G()�y�"�gah��@�{NC�V�1M��AvI,3	M�H��:���:�G{� �<�}��q�(�vW�� ����3~���b;m��ͳ�_�l�3?�D���IܫՈ0�5IH,F�ȃz�F���A=��nL�l���:�:�)��1y�`.��U�ךf�wX�0�Rt��s1�=n͙��^�$�#&�Ү'ɾ�kdN~�#8�6�35�q�*�D�U�+u���Xy�w+V��!䚩k�.c%x5a�>}��xy�GJT~��������H5k����(*��)���;�t���A���2!;dR
 ��z¹_��!�Z�1�-�J>0ɪB�c2j���C�D���::ʞr[����3|p1a�������jE	��|���¤��~&��alRZLGw���\���ʠ#E�����8М�Z��6
�����5��f��|�F�P�=L��D���"�)�����������{v�,�w^ܵ{�sb��b�.�`��S�Ah/�ZJ}ݹI:�k_0���ϳA��#�x��*í������j+G��~�`�6۪���qз��:$�Ȕ!�q��}�Y>���3Z�3Fb�l���fG�l��Hҽ5j�kL�@�x�^nH��z���l~��>�h��s���s����@M���I{�3��a��li5��%�E�}�9��<��*LϿ�h<�d�w؝����o�&& �����9�/P�����&�~��=n{�A��`��4}}ҕ"�j�^�Y�y��A���Gn
���ý�����'�V�~i\1�Im~Ps,����_B�:#M��=!�SZ�:�|8�#�Ʋ�p���BH~_mw�+�N�O,�m�ւ`�n��\Ahܧ.���yqo r��]��`'lJ+n�ݩk�~r�����9C=��`X~�r$����m��Vg�}/C�h="�6�`�g5������b�t	N� Aɉ��B��*����K�9@��7���5��ϙr���DTࣧ���*1�$+o�P�fY��0V3�M���o�18̅���|��hPY���6Cb4������&-��Fb�jY+1���r-��?�J6t�b����5o�p�5������%#S�ټ��-�7�7��tU����Z��d��OƸX�r�p]�[��~}�B���?����K3�4�J���^I���RJ@��?g��0/���n�>&D�M@�M\�\��y�Fَ�T����`R��y:�MN��jJ�؍���|�,�k�y��b
�#c5d!���di��j]z�PN]���5.$������E��	Z"��ڳ;��߹P0weJS�G%�9|
�N�Z����X"�떚�t�c��l����N�͸�@[[Ly� d).�)����Dv������bj���b�ۚ���."��#��i���|�VYBi�4@�E���}0�}u~��:��6�lHa��$�K����]�W���M���� +�flKϼ�	!��
��?�3�o��k�2����Uo�~��0�-.�af����{I�������T.��=�����(!vB	�����H��(����O3�&_�r|�
K��i�jCj�\� ���H��p��xR?���q۰���Y�Bs���n��
24�_}��b������XS�9�c:�Ϗ��I_p8�����[sQ�h�}���i`����M�2֣�;�o���yM�(D�F��gv�D�Շ������硛�M���o��p~V���%�&O)�"�q��?��M��J�2�ڈ8�z�,e���H�@����h�=�@��e��_uu�|7z���@IP�� %O'08�,	5��9F\a���@_	�dGS&�^�E�r��@'�����is��<p4nMf(�Dtv�PIZ�R��s��Ʋ�&�Oj�MW^,��r���[c�3�9Нe�l'q��^s~��n�B^h;%�R�t��NA�)=�= A�D&n amӆ�j�X���O�?�=���u||i��l'�&Jb�e�����r�l��Կ~�'nHƕ.mb���R��6�N�&k�V�em��-�D����W%2 L��mC�"Y�"a��'w�Mr�P}�2tr^���A݆<1�I佦@��2T�>t�z�=`)���?]E�g[�k��h�S)��^���
�Ԙ�L�
r������N��E����܉�żS2�W�<H{f�A�	����s�I�-ZA�$��t�y��"�P�)а��֫��f�D��^�C�<��j]��7�eJ�U���(��Z��"�JU����Pgdh�
<Y<3d��-����2��}պAR"i�u��HcM��"c���/�ii�s3�b�VvP`K:$�}M����$�5�G�,V�9kjǾ����ԡ��Ԧ��l�=I&g@=�U�q*nlE�K�Idz����g�B�-{�G�$�=����G����3�|eގC2�	��<朳BV���RӘY��6�I@��5Pw��l�����Rټ\Va%��1���d�����&��A?���L���-�0��.c"U| (�ru(z�2b8�����{e��P���x��+�|�AС��'���/�D����xiO���*�K�4$`�q^��M3s��;�P��U�+��!H��PЎ��?�l /���"wh��ۧ�2;Nz������C��
��s�V^y\�[��(�n�j�/��/N/E�M���������f��A��0��<���C� ��T���@��]�DK�OzE��
�(ѿ"�U�B�=����}����t[Ē��F�E-�f4���V��t�6hj+%ai����m>֗CH[�宛k�J16�5��O`?s��-I��P���r9��;&����(�xX�P�V�[hj<���"�¥F����k�A��։}h`:�M���O/�"��N���w	i����(��PR�9	=u"����� ��ka����B?����C��JL�d8����(_[����`�gyج���8��~��[���H���P�U =ь��W�__ʽTnCɼN ����>�H˙�\�� �/cIH�&4g:b��st`�_��󨩪�����nɱu�!�Y�:nV2e$/����:G����k�OW5���>��bo�B�+��Qv���v����ș :�Mo�z�%��p:��K�k���鳁���[����.x~.�{�����
��LO���[}V��
5*Iu8g��̑�O��.uF�Rt���!�M��:�2�O�?�,Veo��o3��s�4V�2�`��O;��^��Ŕ)���$_2�&�о�M²U�P���h�����ƒ/����\)���*��y���y�	4�5�,�L��&��) �7�`��H��z~����HBT��պA�;�hL�1Xb����T���W\�:��L|��:eРHإ)��Fd)(=$��BшH��/���o�nӇ��4<�{R2ӯ��A�\MԴ�����GT��ăn;�x��X%���)Y���i���dL���r�v�<��v�Sh�����R����p��
�Ş&�$�/�a�s���w�NJ����3d���m�q���*�1�+�}m��B;7QV��b&��j���lu�y�+�c��  ���O��ifA�["p�gqZb�i��UN|s��C�{�yB�H��`�T�����N�YH@���J���<�E>ؙ5h3=��b ��CF,N�5M;�8�F�>�B#p��@�pgt����-�Zq��k�6om�Itc��v6���4肁�غ�!{�?����:"�r��B����R���s�L1�EϦ��S�=����1����{����g(����;�_BK;�WdFR\����έ��!���������tZd��6A���˔�ׂ�t�]���Yd��9��^�������-����^��'2d���^���L��v���J�z��'%pՊ,��iq̠�:��B��~K�l�n�r7Jh�w��pA3����lA�E�	Z��Cg,&L~� �}ԗ��_���i˻��u���~�+��6�ؤ�J"�':��Ɏ���<E�C��D |�BCVI��D,���Qց���R�%����MI�q��!,P�pKu�_��D���9�r�8�B�c�ʫ?�g�f�o����/x�D�_�5n�P2�sp�a��ד:�sA6��Y�3kmɋ���
����H�u�n/�t�%�Z#��X�R�(��M�P1���!@T�xk�(8U����"L����mSCL��R������l���[����9C,/���6 yM����5A(����4#`M~����w�n��i�����/�����/~��mIpػ3P�ƴf���ZREv�S���&e?
�,-F��u�)�w��� ϮQ��?�C�.B<LS��ф@�o�{Q.����HCx����s�?Z�x�Rt~�����ܶ�%���凧�0����j�����[�9�ld݀���2˸#�c|+n��n�qG���R�|���͏>G%��9���Ҷ3,�c��_��I@}L�r�0�-T���G����1�:g灓��fT�Ƿ��N��dUa759ds�;K��r��]^�U홎v���`b��/4]�Z���q�p7G�������v��oY�C�4����i�`3ׇ��a��)��Bu3�xQ�T�9ʦ\X�J3��Wڨ��G���B��=���p�v�ȡj�w�Z{T�b'��R#X����mŠȫ�EJ���S�Ih��tb�~��(J,�� C>9^̢ -{��5��4	��-���cb����L��Z��0h
tNM~b>��ի���u��|!В��1w��b;�*�O��Z�o�3�i�@-��b�pm݄�KJ�%)�	��ˈ�8��,t�������Z�m��=e��O�E� �S�3��g���/-��$� g�������ǣ��&���J�F"q1���P��?tq�b���=}�n{ГS�q�M g�i���v���JZ�.#/��
��"��6�,Y`�~d��Y���-ZE}�F��>�.I`��
��&�����.U�<%0�o���R�o�T���5ٝ�6~`����'��!<��6�UɛH���%����`g��"<�1�zl�[�toz�@�MI�hS�����Ԅ��Y�l1C���W�������r���Е��A�S�YP'{�e\�)��(W�N�sG���eXAv�HV�� ����og�P�Ǡ鴹�-ːd�n���d�͓֭�_(�%WԔ� �+�ׄ�R�Ӯ�sd�j�C�٬ﯱ�^q<+Vd��:�������f��q䱪�s3B�AP?��=�@���!����P�-�����P}s���	�/�YSѷ�-����_i�[����a<�I.ō����-��i���;�<ī����
6�Sv�z�F�mE'��/7��Z2m�:�wW�GXU$6?<�=�m��e� ��E���'f"�Cj��oS;y���@�/l5:౧���?�_���
:��=��as�t�(�	�8$�#�����6CmY��3~>���mv��6��Q�ou�đ_��ԃ��e�0����6�dBҗͺ��;���#�A��9�ݓ8@n/���z�cau�����Om����)~�D6*�N�Ǖ�+x.>���K�'������+�I�Bnm�z��_
j29ׁ������.������3 �.:��pVpV9Dn'�:�?���
5t\ē
5t�
�����Y.R8�?�� �y�X>p�QV�朠a^�S��\���J��� /�����#pA���`�6{sL7��|�E5���Ib�`��ލ���E/�DM���-R�h93q#�Xw���go���qXJ�g�"�-Ԃ��܁��eK�?���݂��a1�=9���x⻥�;��vۂu-��9\s�R��v�����@�r���Ix!90_��Ğ���s7�O\�CS2��ʨ�'��0�K�������4�8������'�;{iY�Z�I���JEl=R��_r����
/ƊO�-#�C����2��%�I�*R-۔����b��Ĵ&ۼ�`���/�ݚ��`�Y�로��PM���dU��7�`���n\L��n�h��O��X��:8�}y�\��)7{E��e~��(��D����Ppɕ�G��4	�%V�0�4��:�d�˫�WJVF��cXg�@�Q�R�gn����s.ʷv�|��z|W�6�'�*1^�SӦA9��@&u����vr8�*���Th<'�30������� ��3��(p�ƕ�&��XD�\����7+M:5���q3~�΢5�%��Z���0-��b�o�������u��t���h�'���B����tԊ�����
g���A�[�����V8÷���B�C�q�}��C� ��
I���(}wwy�H��	����?�;�0����-�G�5f}��W��q���L_�Mʺ����a�R��S�ι)�[N�Sb~_��ҙLyو� � ��"�U�����r�#t5��MVYK�F�.ӿ#��g�Ʉ��b�6p��"?c�`*��6�r�{�͇?!��0mŌ6T�zO��vxW�A���<9����:]��f4�d�~��0m(y��j��)��5�L"�/��y^ĝ����Pz���E�?*�Q�k(�~�=>�WLi��:r���P]��+�����8 �S����/=p���'��v�٣H�?�e�eF(���,}@��,�rv�]JH�n�c��Jw���D��B�2�U� �[S`��=Z�G>��lz�6��bm��&'�˪�%�y��)`�����b'~�&�n��9��ʧ�;�YLxJ��'ޗ�>].*�L��=�)cĿ��� �.:1�}�����R����i��u���g}nkS�Lk��n -�!�=��L������m����;�瀹z|�j�T�C���%!?qu�=e	�˻2��/0~��nD��6�d����FN�8�!���e,{�ʲ�	�'�?�-�?�n&N��,/Jr2G��OCG`;���>q&�Ǚ��BQ�Sl�ޅ0��ex@q�N$?��OUWyJCj�K�袀����#�1��Qf�~-ca�Zm���t�lc�)����[G���}b�S��J��O�{���`���U������`mS\}�'����V�T(RKׂ��4�B9����J����"��8bh[Vé1��\PD�
��F(��1���Y�Y%&f�44��.ta�⋏	P6
�184�c?�� �4I�����pL��.��^��R��)�.���#�8j�Y�f�(�禯|�q:���)9���t
W��m�o	Tdo�����O��9�{�a�˿�$Թs-r�\E��$�no�C����0����I���m��q= p��Um:#n=	�,���0-v���_��� ��s�צ�N)ZWq��&e	��
I��x�J�Ͻ��9�S�.CQ}�P%N�t��_�BLH�qӔ��0�>)K�k_Ȣ�!����wdF�w��� ��:��|��/�7h<$��>;��\��3�#� �*筓A
�j0����]���#��(�ա��ڟ���Q!w=}�_7��o��u�y�M�u�Blܰ|��i�����N�H�g�_�� '��"�SQz�@u����(�UD��߁?]�3���p/ C��$D���@�pB�w|�;v&�,ɲ�%���eb�o�^[���Ru�=ǉ�!t|Co~fhG��Y,��dzR")Yh�G	i��G�<�`���1�/�C>���o���jaO,C�C�0�ur?Ω��q�#m)�FeA��'�o��Y�R��G͙�E�5Ks"����6T|�wn"�"H�u��Y]H�=�2p��Ey��e�F� q N�NDE��e�s�ⴖ�7a2x=�/�)�4�-�=?£e8I�Շ.����t��F�L�A3Zq�.5W��t�M5'�JCcg���Kp��i��=�S'��>�rkȂ�nڦ�5��\�Q_���\����^!! �g�|(ud��؂SB�+r�~�g����36.�5���b���]s
_P�2�RӐ��!�+���ӫ?�F�r:��Z7��S�<��v�$��S�[x:!<q���H��Y5P?
|�}�[�^<b�aZ�XåJvX|h����E(�lĉPu���h����U����>�]��k�ǎY<�ު#����ϯ�`��3Pm��֌���*�?Ɣ5��t�s�6�S��s7`7	2%3�V�MDm�i����������|�x�;H��
J�(�q�cN�5/�o��V�������)��O���FX���0���zN_�E�n����y)�#�EP/�5s ���sn�OI���Yv���q���c�AQ�oy�yYs{��� �
:`\�G�e��Cl���X�F3�����M���j��w<2��^�,�O�`T�ɇ��	�xe�3�?<):g��u*�j��h����Z���� ��L sg�iWaҗ�8� ��8���؟?�V� l�Vbqx(2�,�J������&w-yy�i�F+]�i�1Xo<*oT;��_0Tkk��X-�W����-���r���%p�v㐾��WkB����i��XH|�,;�����*ǋ:�1̖{��!�E��\o	��Č�7Q��{�t4
=�����[�YL���EX�ސ��%�V祢�&i���n�VL£����&0 Ф�����e'���;N�*(���a�v�ɒ]�v�4�˼�MU�Ϯ�w��N5 ��v}��}'�PS��T���#��P��1Cu��^�1�"��!dS'h�g��Vy\��	�� MM[��M����潵�J��K��'u��1o��g����ܗ�}x��7.R�R��U���sDL��_����N�yn�}K8L�Wޕ��������DRl�<38Ѯu�㋌�0�p�Q�B����Q��w͊�9��+�8�'5z���v�
kĨA)�}�ϼ3�F�Mq�ԕ�㼝k�$Q��8`� ֒�4ۛ,��+'�;ݨ���E�'SJ�ѯ���AW��C�wR�l�Cs���`�9� �%��]�k0573�5S�
	�W��D�n��2=3�^��uM�_3��x��Ѹ@�)kE5�,�%�ś����g`k{�Z;�J�� � y��[T狝E\U,jwV[��m3 ļ�Ы�~o7G/��������Ĺg��wޘ�ڣL쀽��e��R_$�	�2���ę>7@�f2�� iL�D�v�Q��s��|�>�#���H2F�A��YүX���Z�O? ��ب�lU��b�Y^�At��5����b0M�8h���ZE��H��w�u�\>�1��c�/�GN�ۦ�r�@j
�k?W��{H�1��JP
�d�� 1��؏�+���6%�{$���w[e�8��tťE�UT,�N?���X�y��&�kQڗ��(�ey�2���nf� ��^PTꪏ�͊+4Y>�`&�!���f��$�A}����44̴5uS�9��rj-KU��Ñ�L�F�[pZ7Њ0��5«�m"�E��~D�G�sޟ?Au|g���P7=�zr�5�
�|�w�ŗX�;v�$f�������:A��F��D��D������p���S���р�^Ў��?��UB�L�&��O�>*�>�mکy,j��F�O�n�cRAHe��*��&��L�B��n>�r�J�<C2���� ��]HD�Vf��=f��u�\���.X�2)�?R�_ǥ��~�o�_�@���!v?�M�Q����{���i�ꉍ��DK�4�`����ĂˣO1�w�X�2#e�50�pr���ŷi���o�.A� � vY���wdC_�n����b���S;Uㅬ8J�>����F���F�A)����Q=Sp�@�F���N3��X�r�T�P�x넮�E4#S����.~A��pj�q*�������b�D�8׫ڗa%w�8�-a�8��#cymQ�lyy>��1�Xmҕ]M������-�z8��r�!�2:׋]t�UDx��"4!$n�\�vz�:]�f�Ɗa��0}�4X�]�|����V_�v����-��&�����ګ�UE�n�޲�n��t'��)cS��Ed��8�}�K�J-P+' Wsy�ijJ�f�6�MWJ������Y������N��WB�m��91��]��<
zf���������p�=$G�|�%�{����$�:9ƈ���%�����`:�1;��� �9{�I$�G3zi"�/� 9��R�Od�DУ~@��Cg��e���0���������U���~o�?����"�;!$�c����f��d^��bbWց㇞(�\���SM�H�w�uJn��`�9i�[�ƻ
2`�$%p�C��we����;�/LUe��h��j�u���!���jp�;rpQV����n�O]�u�s����f��1DO��K�����|Ҩ̽+{v�!��4y���U�%����Stڷ�llqi���OE��Bԉ��\#�'t1�o�g53\\</��5t�1�5�;���5�H�̇���,��Yz��:��Cy�[Z6/k�5�yO;�]�ȨK�ߊ0%~�����l2�+���$)�$|+(~�h\$Oꢜ�W2-�6SH������aO�����r[�wI��\k�&����:����/0��OFo��4Չ��rE+���X�����Qo��ֹqQ*�-Bײ�j��gA}��D�{kE������$=���na!�:{�d. ��H\��1rq�!�!��6�`��M
���x������ց�^�&ȍ&MQ;�kۉ��l������d�
V��_���� ��H����UL�̴)5�<�������mv*�uX�mIz�N�/� h�e2e����/�]�����w�#�H">�o<=-!k&5Vƽ����i�-�S^>��R��b}����VnɎ@�kw$�����ۃ�o�����&���Rv�;q�����3���P���-�����,��7�����z�KD5 -J!�3S��B/!�-6���Jې�hO�E����|[�Ҙw�ǐ�����Ww���V(�)���O/����EU�c��<�"[��]e�?�X��c�o-X�C۴��Ȭ(�z�n*m�5p-HyM���kQ����>��9���J'��T
Z�K[*h,��H
m�>߯f�`
Ĥ�J�����	�!%:S)�h-�6��Kº:)/��*�ͅd�Ÿ6M�ҵ��~%�*y[��L�/a��W��ט��!N�<���N���X;�b��e~nq��m|lf
�x���=�ղ���Q���)�7��R�H�-;�F/5`l͝�5tˬt�7��_�6���mSq�o�����L
d/�0�7F+�J�@�z+m *�G�%����A�m4+�l�2N����̡�8����
N��p*����3�?�It[Ƭ]��M�eS*oh!�������(�f,ӥ�#�;��ݳhŇ�����=�
y����`Xw'y E�ť��R�lDY_��@���jt���Bz�N�ݛ)Hik�	9EYQzƝ
H�Ŀ����j`a-	B�-��ź��Fd��J�9'}��
,�1�J8-�/1a���s�$P"�A=�"�Of0biN Dj$�2��6������t��[Tz�O��K�B�`��P,�b�ٜJ$�R�a[C����ͤUt��:7LN�b�t��K�������?����ԝ���iuT�`w��4@@Zp�~��)�U[�~pBbݵ&{@����jᓖ��̇�R����I51���e���?�t���C����R��:l|Y�u}R
D:1�8�s`�j H@�{� �����t�"Jȝ�E��Ιo�Q_klDTf�xv��D�$l�x�I��D4�V��MG���?7�<%
w0<�1U艘*hN<B�w��^2|�KZFMvL�Q�[р����1��B��XI�K�ژg)���A�D��.��������ԧ�$1e\C��;�~eXϬLtt�'���~�l��vy9ܓ��X!'a�m�hCm !l��e.�ӆ���D	���̱Qzl��v�#�o̃.��$�DB�/�Q�Fc�D��~�o6z��a=�e2'��<�6�@���)E��Y�3*�NN��)�,��O\�I(�?�(= >�Kg����/��ጩ�T�#��E����f�ʼ�#����8��GFXoa���٨����������"��q#�'���j^Y:g�j�<�A�C2#e"��Q�]�>��%?8&[� �(�;s�|��ё�~V��R-��_�:c�P���x����^���7�)�*�G�2[��@'$��:�)MH�~��칚�#��D�����̡��IR�m\ZP�:G/���|T�7oa�IHx?+ы��V9~	�OZ3� �F�f[�2�`���[!���܇�[���s�j���}^�oF���@&���Ϟ�F1E�!��|���*�g&Ȭƭ�n��9�{Xc��ty���~vdc�琬����c�4��E����$�:����l�y]�0�x���<�!a(��]���nd�R�|�P�پd^;�� S�%xs���tH��踣9#�̻���9�J,d�Ԁ�y�|/��Y��tNt!V�#���9�$j��+���<M��Oad�j[��<n����f�Df�u��a�S�- �6�O�l���=����(\G�w��@�X��c�񼌌�ṎF��
	2�*X<�����p<'��"'+�إЗi`�w�Hvg[$�b�Br4���R�e��9 &����%��%i��1��͂�:LP��C���� �j��8+C����.�,G�hvp*������'?�5����@�E��S� BwO;7#�$���~D�yyc�A�g��|�����ڵ(����\n9œg��m��b�g`c1^*LC���٘�5���`���Ú�GݤH�m�9_���ץ�; R!��r�
_r�n\�--��^ ��9ty��ř9@՚�Uɓ���{B��vDU,�����1�}X/��uA-�#���O��f�X!a��	1b��>�{����-A_�ɡx��?d��N��V���P�����8d}k�OY�,VUhnҤ;o�y.G�_@��nwVT��C��Rb.�A<u=�Z�\���y��E�sZ�����4 4��9hY�<�u��1���o����R��昡���+�v-s^�MQ����� ��y�2�a����c���\Q%�xp�%�`y~-�VV�Η�y�
�)쁖��08c�>� "�M�=Y����4�!B��{��l��T�)���o��I���=l��]��~� )�&Y��5s��/�:�,oq�E�ٖ��I�e��Ϗ�h�`;�fLk뉋Ba�T�K�;�2�$<V
�ԸҔ��SF}�f��+ٳ�4��GFUU�[^[�~��Qt��sgf(W���d5q��I���D�WR1�b�:���uR|�Q��|�b���m���䢔�Ev�#��.�myJq�X�@�gf�����J�<�=��3V��0�{-��W�ܑg��waF� ��.�s ہ�@��8��ADE1��F��ը��w=ɩv�N�t�"<O�X�a��~�D,<ޜ���L�@�q�k���s����D_��ʝ����] T6�8,b���^��J�$XP�!���FCtu����Ve��~������_��قFnc�zhX���QPG���"�b�Y�7
>�a����2��T"��
 mA輝�>��xb���g狮���쵔�<��
+�n8�6���m2㇊Li�)v?��$=C0f�W�*g��;C 3Q]i�����\!(���I,�����di�D�-�/3t5HDc�ׂڴVδ���#os��p8D�9��@����d ݽ���H?q��ԛ]�.�$O��[D2�sl��	iT��ᇂv� ��O�)��s��h�;�FD��ʾ�D�5�����92Ե&�E9�ھ�~��j�a�sN��4�U�a#�٧��M�3�/��t)V!���"�Qo�߶]�@KTRu,,	�_7K�~��!���:_^Ȯf��>����8"�L�i'e����'��0)\�=���א҈M딅����C�#U�!��z��V̑J���s��Fiʵ:��i3��/�nu��G���`��J<q�3���	�|{����o� 2�a����>�B�*OL�����y?�J8�&����=�j|@��=���jHXa�g	>Z���g��(�R�p�C�s]J�p1�.h��%�0��d��x�rB�M��}�t\u=�c��{wa��Ǧ�@�i��{��#@/�����f[+���⍰`wM?M����!mj�3C?Y�_�n�r� }U����T��qj���w31Ӳ�:J-о3¡X?�v\)u���(P��n�t�^�ߘb5�1��!:�2�юz��ߟr��Aw8�X.&�<'7�Mq�>����G~0��5�;e~�'��%; ���_SW��]%_�JC��Y^�=��:-�}���/+&`^�(� �W�d�b��A[x�JE7����4�_��\}bDh���/���;���<1����(��9��h�v�]X�=vt�klΙ�b�ʷ�N�cl��:S����<�֣�bF"G�v��� ��ˢf�PD ɭߋ��z��|[�����qZ-j�I������J�[��Lͨ�TJ��F��as��<ߞ�j�gџQ�[:I�"SB��ks���8Ď*F��\;O��%0Mo�a����g-��Y���t8�c|�ӟ�س�
��~S��ؕ�6k�ě��U}\�o�m�IW��zU�az��}	r]�,gۿ���2l�m#�q��l:�S��`�u5�?���="��c~��\6��.* �^�v^{;�5phm�_��Vz,������ �
R:C����sCI��^��Ek0�-O�oĦ�s�N8�7=�?�G[��o�u�]Nk5��E�������iqFU���4�����좗���"<@H?�=*�8 c�6f@nM����'�[X/)��AF�T/G��K,I'�6��؆ R~�xB7SY��6Y�׳�������H�&����!��Yo-���F ��l��@x�!���ԙ��ȫ��ܳ�b�IwA���<����&a�z�����j�Gd�Y9��D$�*�����(�z$�<�:!�&�ψ���Y��v��P�BkR��(i����>Je@X0��gQ(�ļ$ a*�������Z�q:�������S�=�Q3r��)�,@􌙎�/I	hV#9�|qD�K��E��\}�`��I�z�����݅��GmKQ�$Ib�]ˎ�C�?oڊ�D��b�HK��x���_���\��R�
#�s�S����bv//T(��+���B����/�����ǩ�נX���$8��퇀z�KJ��aY_;�<�.�S��B{/��5{by}����x���r#�y�䆘٨���h�ff�8�������3�k�Jt�>�B�om��(J.\��ԝ#���(��$�wg�ٜ���{���y�ҽ��+j�+	�~��_�ϟ&��"���cVʹ�s6���p��"kf����j����~����`;Q-  `�%����l�����Z�c�������m����w"��r,1�tV_��`�;"��%ncl!hؿ�s���:�7���N�7����[���
=Pt�=ʂ���O��Id�S{U��H�!����+��o(`�$��=���s;z��Phs�ܧJկ�C�+�(ժ�A���r�/�����$��J2���Vk�鈟�Qr�W�Z������O�E����3�T�C��2��>s����Lq�[r�
z��I��k�GO�?��;�<L�Mx�k�U@7߰E˱,F�-o���_�������*Wi���u!�@,X�i�Y)��1�`�b�K�L�ç�|�=��Q� hg�f�n��s-���W�� �L��:�r��ls�o��hL�uZj�����SW,��g��r+�3�f�6p�4S�.&֓�#��Te���}�O����mD��G�e�����1��C��n�b`-j�э�7�km��7�Ɩ�.�۾U9��`�S!.�Y��41����@�9JJ���M�q��\U�YG��o1�+1A#(���l6ݴ��S��z����ޔz<ɀ.Zɪ	�մ/���`nfc�V�)�\����Mv���/�P�٣ �W���M���Ytl����/-ʱ�h]m=6N�A=�Z)vZ` ҕ��?���z`���gU�T̋ߑ�%Q�׻dĵ<������M�	����c� a�zՉU~�T?g�I��({~\�Q4 1(0��|+/_���7���#
t���0��"d��B��$/���gs_R<�g����2�^ߓ�PJ��wl\���{�[vE,��H޽5/st ��9Uh���7�&��#�I�vp�Y�v�ʹ9�R(l�c��uN�T'g�� YaR�;Xٸo��|!�_o"�@���/T��(���ν����`s-9L^wC;��t
BG�e��!��/�  'M�Su�I�8{�s��$W	2:�f�K�YM#�l�C�¸|KRp�3����1�{^i\SC��^(t�4)$"?w��gxJ'r�˩u�6�����L*b[q)��r�!nSY�����f&�O���:�6�l��C�dan�^�M�ǈ/��9�-=�7I���"Ŵ��3t��1�삿�Hy�+#Ș������-m���Ax4M"��hw������|�B8�����	�Le�1�$�C��j�W�_��q�<�Jp!Jp�4��ignM =M�G����Ѯ��p1e�j�P`�}��M,IN�_F�n��zbs{��[�Ej�5j��?�>Q1�b��1B�9�$�E���6����M�T:�yfKF��p���C)"��1�k������4-ʔlv$,H�R`��t*�Ac ş��>��%Nu�����S�s���e��ɀ3pw������{���xj0f��I����s@���4��0����i<2�}#�0���z�-��	��)c��g��6ܴ�!" HFD�=���R�%̪�"��*�Ԕ�))�?k7Y�ZY�J�ё���_J�x���ƺ���������Ӑ����!�}~��b��V��3�x�˟/�#K�Gx�[��Gbwv��"J9�: �J����M�٦�v^����_)������"_��S��q`0Nm��xA@���H%�/{B �t�҄���������$a�!�
�ɔ�ר!Ŗ����$�M��lפ���L�"���m�V��?A1wf��R>x�����|�[�r��$�*��/n��m��+{���M��v�����^|�6�Bm���W�5���-N�f2Q�$�����O�'@� �H��8����ݪ���y�:�$�:R��J}��e�R��k4A}�0����/�<TBű_�&�,��l5�{yAը�3�Rob&q~�̣s]�����*��N��s�L��3�]��%dަdt���>�r �0���j���'m(:�mTy��S.���z:�\��%��U���`6#�p��!�}��Pʠ�����bUG_�[@���ݔ?s�9Dͭ�S�
�.������.x�kW[lw��=s������{B�ͦҍ�-�Y��{`f�.sG��c���9P�o�0Х��F�5��ݹݒ���X��E���8��r7u{��@��CcS�W �
�+�в=�d��MO%Ohݍ�A(>-����-�1�a@ �����1��2uj�"�9����H�Pv\��1B����N���-������`M�Fn�1��Μ]��~��~��[,s0�ןh�v��Ƌ<��Xv�G�J���x2�2��^Q��b��W+L:� �2�����,��@���킔��m<�&�*�?��K����dz���=�#T����c���]�ۺ`�k�7Řׅ�~z��{P�]&�L�Z�tE兜\���3���"Y<��~�4����=�n� `ki$�'��6d�}����M�W@Ov\���3�n�޼i+�v8	�x��4�U�j�&�b�Կ�l���Ʀ&����X`�5u:r&�\�qO�����6h��ԭ��}�'��M#z���[K�sW!A䛻�1��N�o@�Tf�l��8N�פ��V%J�۝Qߵ,�i`�Ć�ӯ�U�&-D�0��o27�0K^�2�������-M����qu��TY��_a�[v)ͤ��,�88k�����CS�F����)��,�:�)�*�.��ne��X .��ˆ��-Ch�B�Q�����T��O�}��k픶���N�-��o%F��-�'���WIf?58Kգ��F��Tү�zNSwCk�9?!ĺ�,�2�	��� `������E`���b�E0F�v����[�gHn�l�t	J���F�YD�[ei:�!��Iv5�ň��IJ��(�BnD�*ߑH޼]B#N�zҤ�`�f����j���o�������"	�rއ�&!/����W���׬TSS:�ITZ�<9����7��,���e�]�S��a�l�C`�ԑ9��יlk��4vz,�i�f�i��2�m�aW&U��p�Y[mb���m{N�}�H�U0������T����W7�G�|�%�Y�fRZ�����~GD�;R� ��b����f����bÇV�\�.#�]p����Wʪ=h�T6�X`h ���Y���<�������=�6,v��������)�t0�,��L��l�J�{�#E����R���b.is3�̢���;�w���Z*[��+�T$Fii���Q��x_㨓-�-��I[��2i����W���lq,���2���Ta�fi��@Y���19.�zi��iF��s@8?�9j��iT�ذS�\0��z2]�^S5�ݷ����	���=���0�n�����H��,�-O��X��D�m���-uz-H}���3ݳG�sɈ�	}��o��]c���Apð��ŕ�����	�8�x࿌.#ˡ�ĭC[P�(� �&g�g��ż�m��A�Q�f��7��7�4cxR��TS� d�����~�Q��,)c�?%c��%��d�^њ�JB�9�;�k[d4������o��'J�n�i�[skt�6֯�|�R���sS�y)��gXA����ΜY�
��P]�g�lr��$YB�1�c�I�� ���)w�D�fƩG��L�V)iJm~�5�?����͕�_�v1�/��9_��x0�&��Oh�I@ �ft���ť>���ȇ/����_��)|�L�T����Bw����������/,#��y��ʚ>_{c��2�[��E{�gP�������-���Q@�ǃ�+�02u~01:a4{�����̦*4�k�3`�v�o*���):���B C�{���~p��Ȯ	�G�}�P�Z�X�~��k�6w�8CҔS�פu��r�k���*t�T�z�QL��º��5ۍgJʎ[�&?5p����I4���R��'���7�jGpv�^m�+�t�g��n��v�84�W��E�#�����r����g"!}[��,L�+v����xJ�sZ��)���H
I�|����۶�b����	�	؆N���X)�(}̮p���d_#AW�{��A�hC�'�?+@��S>ѵ��X��t�ٿ���R���=2����a�$<1r�N��(r!�@�kժ��k���6i�?�%}��[t.��;d�'�3M��nw��'��E�6ԹH�ґ�PC$��T����ԓ��ל���jπ$J��`B��9
s+��Ѯ��Xz�E���T`#˝�ӗC�z�(~�v���X�5�O�Ă�Z*���0�
��lL&��~9O|1��*c7�ĭ׸�m�X@~~��=5H�w`Zg|ݝ�3���^d�Hb��/�	���_�}�}lr6��-��^�t�V��~���o�a�!��NŨm�+/��}�[�|���+�r�"X]�������l�;�}�s���m`/x�Z/[=��XT�3�~�W��'�W\I�	,�|T���g��?,�΂v����{	O�����پ��[ ��z^��'R�y���AP��Wjh��@�������e*�&�s���z�HF���rp����W�e_��wL�@�]8 ,����-�t���QWbGG)��9a{�]����e�hF���5~�_�]�r���L��T��O*�7�oT
x^M .�S�!dc�_11�ʜT�M��X�c�_��VT/c�p5M��3r�۶��Z�}4E�6�Wד]�T�ˊ�3h��3�=���%�T�4jT�}A���G�O���j7m	h9�x��WIn��ƴy
y�8a�F�8㙩�z#O}�/��G�h��AWE�l=>z��L9�I�Xͣ���#��<�+A?����B��]ai:+5�,����,���z�"���1��Y�ΰ��uV���f�����O]�F���*���r���w�����0��%w�� �cuw\gf��V�(���O��F蝞�V��1�d ���+mF~x�vY�����G�Q��{�j�f>م�T������0��a*kq4P�H6X�b¦�'ʭ��@��㐯��m��\�Άwww���I����W�g��Q"�	ȑ���Q���l���[՚���î8B���z���؈��; h
��_6LN��w�#��y�]L���Ei	CwX H�I��N��%���궩���	.�IM�D{DS]���~ʇ9x_�Yd�ئ;}� ��x^�OB�AU7�����^�j����J�v�W=g6��<������U�V��8��x*�S8�8B�h��+��\�l��A�ZäI<Pru��nz�3�=O;$bi�!�1����E�U��Ax��w���]��nO����E��C#�aȾ� R��O�}h�ס+������^0��K�u��\Èt�֌z��n�\�R��`ֹОQw�X$�-�	��f�	�Io�A���EeſȞq��E���/�����������3e���vS:�W���3p�p�]��+Ek����8htZa���i�ў��fTVǟ���V���f1@<\̃�~a���&�l����6�B����
���z�#G[6�V��	���ÿ͖��TU$�v��T63܄s'�F�]0�8g��_���\���nw��#S�<B�K�ܑ��������z�2W��e2Pg<���/W@�Tbe[����Ն��E�Z`�Վ�%�\#F�Z�H:�}���қ�Y�\��3���	h�+�'�4�a9#Qɟz08lu�C�9xus�!?܉���3�{=�IbK�E1�iu�ռ����Ï@k�`�6:A�y٫vRƒM� �%f�uR���yN�'�b� 𩓍�� �����W��b�;�T/v9$r���~0��m�O�.U~�'Q�Ť��ZU˹�Gx ņ��nL���A��Ր���|���$!�JvN;_+a�["�W������|�)攩�1�}�������Lѝ�cy�����D���ְ�GZQ}�^t	���	��)h�Ue�y��'o`F{��
/Ż�~ u�'��ZG�8r��o\��~ޯ��~JeX���d�c�n�F	w��e+X3���o&[��D��{�q�����d�mYK��5�@)/��7�[4UM���33����Ϛ����	�F���0�.P'��%Z��yQR��ӗg�]\yI���h
*L;�`<]��d�IƏ���n�b�����0;9��m9��JhEn	�0������o��"_�H��o$$��1�ޠ��j�}��5�b �&?�(��u�Ct�5~)⻓H�nҟ��� 01��f�� l�����oVK}Ny���ʨ�cD+m֢��;>�,}�]�!׶X�)Q�����ZT
�0��p���N��x6'���	��#6��~;R�Ƅ�ǽ\�Z]a���v���7�x/6��������y�!��8�����$}t+z��W�kw�4��J����5�t��B�]����v��A[`ʱ�����>�ny�)@���?��AG�k]�^�	-�Ѵ��MU����w�YIm���俶XjF�U������6̈́W���3(Wҳ��'h�d��V�W���k܀k�c%9�A:�B���0����8e�<�@��۽�&}{$S��])7F���!�0��H��ݪ��&��B��:��&3Q�3  ��
M��\>h�4�/�Ⳳ9���.*!�a�D^����S��8Z@�[��Ƹ��e̏d+�kjJ�-���{'|�4Q`
��~����V�如^��R�M�z(�Km���P��n���7�/}t�Jz��W�Z���{"������[H�-�oZ����C71zV��AA�R�!t���A�UP ��(�B�9 ����t�B�!�Q�nN���8q�k\�!��̲����:D4�緧,��h}$]�����V�
���~��Z�"����8N�p+��A�����3J���QqB�=<���W�mN ����Ր��G|�=`�}E�E!�sD�Q���j5�aK;^-���j�B$���æ�.�6�x�E�����Q�~%��� �p���u�d��e�O����힜�VE։.�bK�����ӥ����m�J-����a4��N�TR������������mWW�Ep*��G�ߗ�zb,R�?W�������U �������<"�|j���n ~���43�f,�.%1F��~2W�;-�ΤR�ܮ�})�?TK�'�INP���x,a�j����`��;&P5Ɣ'�E�Bj�;2�����b����e����{x<<��5�)��ף��?��[o}j_�S�s�<��&L�.�DZ��%�ɠ1�^�|�`��1����*�{0a�^Bc�-6~"��\%����k�>
�����.N�z)f���$mQ.
���$z���uAjR����[^�z�l�6/)XY�����O�Y&�"����C'/a�FY� 9(m��م
v�w�g�},z+N`�d��U-M ):2�I�%9K���y揯,�ԍJOV�@��"�ӈ\�`�xg�}���Y�Q�����<S2W���4Bہ�9*|^?|�����0�b`�B�MB����iP�J^�]���DP�J��N�L
����0(���Mji�\�O�rZ�+ޑd_>���6J!�2�}�p�^/F��Xtf"�B�߄�2ǮqԔ_�)��a�_:�M��/(��7�����،���_0�ɞ����^H9�|����{y�� <���$k��8On �L�Ŕ���;��Щ����S6�]�o��S�N�O��.j	n�#/ |3�#»�C.���J]�F&R�4��!�+�(Hw<P�44�ƶNk���C"�k�Fk����C��9�C������T�#e���>���v�� t�H�B��QK[ÿ��O@0��OY-�r��1�}? 4"���aY�8/*�W��@��E���Jj઱�My�4����|�:� �� ͙����QG2;�1��X�|,^��������j�@���O<,��rA��[���\G �:�0�-&l\i���S���+�}[�t���Ax�����_Tخ�-�׿&����L����y�e�\�\Xo�S3���.�ӧO0*5���D0��L�'�E��&2?+����O�A�+���=�s�_V����Ms���q��%tL5�*.�i��!�.!z@!���\�9�)Pޫ���ʓb���sLa|� L�����zb�@��^R7zj�̝_���N���U�/���@���
�UGJ-f@���ۣ{��X�LgΉ�A`��!ãg�sA�xq�R,OT�`�9��~��T�Dg
�s�ř�Z)M�h�6�e��E,��-�u84�)s�R����`��S�[�65��ߑ9LğLj�u%���]��>��A,�]_ߞ&I�5��qI�Ҽ�2b�XC�81��3V7$��ƌے3}C��4�`�͎�f�Pq`��7'ߋM%���ߢ;��Uɇ�O�j�Fˍ��8s�+$1a3lX�w���l�܎ϛ����W'�C�?�� �Bo�tV�V��|�����oA>��|"�	���_�W*�P�"�a�d���*;���aF`�4�a�:������ķ"\<�!z��`Sb�1>w��Z-7�����GY��;��y��qNi�.�u����9Y}�uD���w_�Ie7��c\V���"(�2��=y��@k��؅f'9�b��G=Z3�"	Ω?JDk!��������D���!ʩ������!^�crq�"��Yu�-]7cM�s�2�=�3���E=��N���|��w
���Yj��0�^=�({絾���͛p&�Q8|��/F��P������q����MyK�\y��3+�&���irt�5�Kl�8m�2r�m�,AP\�'!�/��G�T}jT����P�-��/�+�$���wT|�I��'#�����y��%�r;�X%��T|�)����;��8��P$,�F�(ef����<������-�x�S�y������v�L��'#�k�?�Tȣ�J�x�d�! ��s�y��=�݆Υ��0 ����Mb.{�����:��C���-���_
���''1^|�cD���������U.�*��~EN�s��$�t�`,�x�[��j�x���N��ag�����	����Z��#'�����ҍǡ�� 9UmQ��OV��0Q�M�s���Ry��(p"��x�Z]��^<G���F���ԩZ�/�93>�P�(*���f��g��; ��l���y; �Y�/H��Z�LK�opm�ȁ�)�
l�j/����,�)�/-SP���-8��at��m��PX��^��r1{W���7�MM�c�U	/7�Yv�7����+���d�1� b*>d��f_{��Q�S�����㑆��v�����$�â�&/�M�v�+���!�OO�
Jl�ԣ,����&Y��أ�\�_�6�tNqgb����}����S���X�����QwT)Q𓦗DC�3Ͻ'Ů!��]w0��\{���s�
��g3,�p�j�v�mAH#s�z�^Ӫ��OT�aW�U���������ǯ����=��龓3F���r�s���?��D#q���ɡ/x�jm�y���+G*3&FK}y�L��8o�Q��Q����ݾx@
S"����j��@o��tc��a�nCP���0V����b�F�׵ 7x�l�fc�cjz4�o�g�[��ط2^(L�ڭx/f�=�8��c�#j"g������5C�c�}�jZ/����]�%��W],���C�"�r��0I'�P�	P��Km��X6ݶ�w�o�TZ��^������)��F�zρ����Qb��d����#�K��&$s�ey>�o0H���x����Y0Na�̯rٓ����U@���6��$-xMg����ݖ�"�tf�T�T8�H?0nA�v�SQF����z�)B=��x���K�3��r��ck����q�u"Z��Dr����T*;n�4�����8b�g �	�` ��3��7&.��5�If���������J�l=+���U"sh�"Ok���nD7q��+������7��� �W7&g�tTsr��2nx+ �Ǒ�}�`�q��J��X�@�����H�{���	a�x��p��'�7/�2\N�l�n$�^�QKE�&W����D��?����2ʻ�����>�}�S:w֕u{s�,�x�����z&�>c���G]��]ᬾ鰷��t���<s�)+�Ճ�_$����?�3���ܒ�1�Ÿ�& Q��+Kh��+������Xr��-) ��X[q.4��9���v]
��t�/�;.�D���?@S�7�7�ˑ�@�,�3"e��Z�d��bBGiS�x�B���Vw��K�IT��(�	~;�q���ͭ/p{K�ƈg�<H�%�/�#�>3`q�5�"fz��?��	�Z�Q���Sh%�d��P���r�H�'����N"N���[JX/�!��'{�� ��l�v���*Zfe����ʄ��%����W���X��a'�c�6.��Gy�K	G��AJ8#ܧ�5���?�ng �ʹ���,E�;8�=�dUm�����)U]�Zs�~�#�pBp��E�H2+�Or�fMW��(}����6�}�ޙ���{b�K���K��F�r�[��z��9�M����9>�K��O�LTʀ�p��&�ř�&\n�m��c���z�uM�-2�E/
w�>��M��`�[D>�=9V�U��l���'ё�,7�r�J�Qw���E�\��|��a�$ڃ�~1����pJ��q��00����c�������Nb�2�$s���>  8=+�/=hb��	k�]��cF;��E�h�o�4�(>W(ubJ,4��>�T�z�7�2���$, ��R�uJĴ����¤lG���bh2��.eHF`ڳ�>�M�S{��H�Wo�׸4 �!dP$t�u$I"�JB�s �e�z����g�L5���KNnqѷJ�Cl&����(�r�KƇ�`KN��`t����Ȝ�@P�G]7'ZrϞ�4�� y��;�������� <��qh%�%Ҕ "o��a��*ޕ�D�æI䈟�z��GҜˇn*�+�k�0Oq��lԧg^{�8?���
a�⃾�}{t��� ��C3�X�X:����Э�1J�Ou>�pc���%��'R��=ݒ&X��K���S�8ſ4�n�+C/�`�g��ה��:���WBZ��Ce�=���}���Q|%{-s�i5U  @��
p'�OE
�GT�(�]^��JC����P�� f�bI2'n�N�ِ�I�M���.�]�h��:���C�����e���&�%P4ʄfZ�L���j�SEM+~��2��M鵧�\Zβ��6����})yLAB��J=�>�h<9�=��ݭ:���{��p"�[&��EQ�.�<�trP���v�UfIM�Q��>䮃�`��f�@3�I�~��"{J�>aƬ�4���ea	�q�Qpl���"���E~��g� ��N#��f��،���g�����v�2���Z����fd�"�����+z��~\�c23�*u�����	-���7m�R����~HEֲ����Z�|�#�Zr1��ʨOAoS�!L���L��vy�K�����E!V;$�EEC^�8����fu�eR*��옞%�q�' %��	u3�X_O����L�ݧyB�����)�f�I��/2E��6�g�H�Yqc����vmL[F��=�E���A�ٻ���|%ʓ]��c�\�l�=�����,��F� �Ġ}�ܔ�S�$�Cc�V��e鮡���F��W�zP�˴́��Ϟ���t_(�����;��%��v�+����8`�dӏ��(���'o��>����+�<&��(rzn�����:�/��WG �0:s:C+v���]��f��%��i&O2�zM��:8�����La��� <��=:K���V��z�+'JzP����X��Pw���Z�c3��OQ��q����B/޼�vr�?�r�lH*
��a�I~N��KZ�s�.�V5[bmIyS�&�+�YOл�'?���$QIOg>D"���rE�iȧ3���7�^/������DDq�P�"{OH�+'�òQTQX����X������ܷ�%J��Mpǰ�h�9`!��&��'�n#|c����&G++�ӑ��������L+ܭ%ـ�������J��f�ū܉p��ӯ��Z"em4@�ca�w����ߟW�$��7ȇ����!��0�X��
����^�����d��3���S��n`ɴ���,�mjȸ7 �|ܳ{�Y�����NH�-�ϝ�uO��w�ks�է��u��g�����q$�}�lR\�oE���"��Z�2�o����e��)������9�s���'w{�(���ӵ�kwf��.I��c ����N�6h��c��%�� X�(__�]���e�� �j~J�6��rSL�jXJ�9�^[�Y���;��l��du���cA�9�M�B�]�Yx�)~{���Qc�������G��1&-�G��Z; �xM� �uy��rhNW�i����pN�R$`��~w��8<�}�cE�0��|�J���{\��2�� ћ!��d��FґM񩣣�X���R���$��h�F��N]\�|����O�bXLV�����A0;��?V�0/1�����ƾ[�{�J�^���$-2�(x��{P\P�;���(���.�$PY���!����e����}rkc'K|I��OE-C����I��M0��qm��{�f�'�����Q��@>��+����	Ғ���H'A�݌�Yfʴ�4���Z@�B�32C� =���#��@����]-j/	��/�\�g��m�\ᾃ,�i��;]�{��'�g��e������׏��`����03�kg�cI��E���?�.U�bPǪ��,����Br8]���?�W�jHOI��ő���JE>#Ș��G��K��J�l�!F��]p������#S��0�v*@�,��s�0L��r�os��4k������l�ܵ3ß0c�
Uɠ����y^&���OS��E1�N��13�/��oN�F���S�Z�}���tRN��f�[���(U���5��|�+e	�v�PۨD�V�HsO.P-�|��}���"���o�=���з��L0�D��> [�/�=�v��C4э��0ı�HA퐆в�����܍*��mc6�Q����o8��2��s(o+�B��z�XPke�K|�7Mև}:�N�bii�qWl�9oz�WA��C6����"(i��[�19��'*��v��ܻ�5��3�{�ϊ��]̐yjd�SO��3��=����[z�dxv�DĬG�o�R	� 1�A��ʵb	7��T/!k��ݳ93�^�����Z��XDժ�ɑ��8b��S�c�?[ծ6������Z�l��=JI�6���E�<��)���ypg2ei u2Рi8��`f��O��@>�y�}F�����*B'�M�d��S|ѓ�mǨ� UT�J������pT��j!�tލPW�4(J�%)`�3��#��6D�<�����7�$_�4vOX�TXm�@A%��b�u��,{�Ԓ�}_8����� ���K�htd,7�����Y;������\�`čּg��X�wm��������Z�!�H��{<��E4����s5G��X�:�BL5�'���T�.�}C�;� ���H�æ,�,��׫�.=�R�'��{{^�*b�Fi�MWu�#9�s�MԤ�8$���:��ym��Щ��So�P�Z�LN:\��;i�Ѷk��Ιf�� �s *������3�}��
m�T�m��c\�XY�Y�E��6�b�g�"	���ÀP�̴�3O
"I����ޑ�� %��I�������ё�^Od�0�l��f�埊����QI,���t�t�I��ʜ�;��ݸ<��-qMV7ݰW�{������&!�:�X�~�w#�y�K���`��-�ag���o{����	�F:Բ�.%�i�"88�_ '�y	V��{��?"��=�J�5v�#���w�qK���%��5D��l�!���(I��$>�K�:� �h�`m�Y�ɖY�2��;w_��>��t��O�a�d�1��T�q�d��S�:��Z���7��\;�c�lᬩ�Bo�<AM��TV'���[�D:YJ����V���}��!�|M?[^Ƿ�{_����׏�EX7���-%��� �Td�A�^sd�������Ҷ5�����3,l�9�)�vS]O6j7bT����X����Wb!�I~�	�;o���Hl{�[2���.sD�L�Ц��{Y��:���&��I$��%o��r�]�t�bE1�y�ĜY�Q&�s�7���ZL7&�g u%C�? !#_�	�al��n��̨Lov�% �8b��҅�ĝ�Bm�ySz�(K�0k��p��m�j�ԏP|PƢ��	�H)ˊ��O��)"Eu̼�ǐ��x33���v�gj���қv�}�t�~�/�˩T�cE-b�R�����:S�l�¦}\zawt�kvx�q���F�
޾��dcU�ɒ�b�(��4��G#�����+��/x��&����0ZU�ԧ�ۢݔ���u\ץ����1�"�����T�Xo6��4��L�l. ]�U�/"m�
�� [+@u�Ix6�X�2���XP6��[�R�5Ϗ+��ڗT4r{9_�ʈY���0���ȍ�����@L�ӀÈϻ���,�4M�,�����	g=%��;�{��'�qҟQ۞B�J'�?���Ǎ�m"�̜������8B��x���{�lD�� �����p[�¥�۴-�8����f�x�=1�"I����L]�*����+�>��L���l�g 2��P1Y���	sq����E/���F
�Yp�aKr����ԝ'���J����_��L���e@�a��y���>ɉ��X��a�`?`"(���_I��e$7�j"�}vmm��8�j{�M�fk����������p�I,P�Y�v$R%	WN>�I8��`/�~V�ʰ��ܑ��7�=$"`�ڕ�5C�1HF��/��*
z���/�,�池��т�ၧd�{�M�L��b%����E�7�g�2��Z����u��h�Nؙ|�yil6�'�lV$�E�YY����c�<�����Vy̨IwJ ������l���u@�2��d`�fKCڳR�� }>D)���&.�F�S����x��s�EӸ3�����Ro�)�)�*X��8ubíf�wg�[�2ը�%���<lsC�h�����M����Jz>t2�Z�Bk��<	�l/19Z<F�g/��Z�ڪʲf�S�i��1^hD��y�6L�20�t��^�?��3
M=h#K;Xp��o?��